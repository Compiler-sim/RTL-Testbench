module wo_buffer #(
  parameter D_WL = 24,
  parameter UNITS_NUM = 5
)(
   input [7:0] addr,
   output [UNITS_NUM*D_WL-1:0] w_o
);

wire [D_WL*UNITS_NUM-1:0] w_fix [0:155];
assign w_o = w_fix[addr];
assign w_fix[0]='hfffffbfffe19fff94400003dfffd89;
assign w_fix[1]='hfffe50ffe215ffee4cfffd0900052d;
assign w_fix[2]='hfffbe3ffe015ffe6e100028fffff69;
assign w_fix[3]='hfffd27ffee21ffece0fffe870002aa;
assign w_fix[4]='hfffe6d000bf4fff120fff830ffdfb8;
assign w_fix[5]='hfff8f10030abfff477fff74bfff614;
assign w_fix[6]='hfffa060020c9000c90ffff84000d16;
assign w_fix[7]='h000373001418000b3dfff9460020b8;
assign w_fix[8]='h0003db001009fff74bfff5d200176b;
assign w_fix[9]='h000574fffff9ffee63fff892001c4a;
assign w_fix[10]='h00046bfff6ca000274000256000381;
assign w_fix[11]='h0001a2ffe240001766fffe2fffed7c;
assign w_fix[12]='h0001a9ffeafcfffcabfffd78ffedf1;
assign w_fix[13]='hffff2fffebe9fffb46ffffdcffef06;
assign w_fix[14]='hffffc8ffecc8fff6dafffdd4ffeb37;
assign w_fix[15]='h0002a5fff5e90006dffff799ffd66c;
assign w_fix[16]='h000681fff605fff50afff428ffe46b;
assign w_fix[17]='h0001790000cbfff505fffbc6fff03f;
assign w_fix[18]='hffff46001549ffef84fff4ea001546;
assign w_fix[19]='h0005b500033600029affff5100209d;
assign w_fix[20]='h0003dcfff5bffff290fffc9e00115f;
assign w_fix[21]='hfffe83fffdbaffe568fffba600103a;
assign w_fix[22]='hfffd14fff09cfff7d4fffb9700070b;
assign w_fix[23]='hfff9feffde7b0005e2fffb780001ba;
assign w_fix[24]='hffff14ffd653fff7affffa8b000294;
assign w_fix[25]='hffff9bffe939fff5e7fffdbe000a2e;
assign w_fix[26]='h0001020001da0000a3000636fffdf8;
assign w_fix[27]='hfffae6000d2bfffcd2001129fff40f;
assign w_fix[28]='h000f3d00013bfff360000a70ffe8e8;
assign w_fix[29]='hfff3a6fff965fff18b00103afff8df;
assign w_fix[30]='h00203e0010cdfff9dcffde22ffd6a4;
assign w_fix[31]='h0017cd002038fff58afffc31fff027;
assign w_fix[32]='hfff51a0015cb000c21fff47bfff983;
assign w_fix[33]='h000040001d81fff760000569ffec4f;
assign w_fix[34]='h000515001788fffc4a000a9cffe9bf;
assign w_fix[35]='hfff8f1000ffbffe49500102bffef70;
assign w_fix[36]='hfff89a000ba0ffff1dfffce6ffeefe;
assign w_fix[37]='hfff31400130d000504fff77bfff430;
assign w_fix[38]='hffff34000869000f96000a04fffd21;
assign w_fix[39]='h0004b3000bc7001655000b0600003f;
assign w_fix[40]='hfffc3a000cc1000c77000f52fffe37;
assign w_fix[41]='hfffab0000bfbffff5b0007e4ffe806;
assign w_fix[42]='hffff5800057affe9c00002e9ffebba;
assign w_fix[43]='h0003b30016f30002acfff58dfff3f1;
assign w_fix[44]='hffee270007b2fff762fff3f5fff036;
assign w_fix[45]='hfff8e40009d80000c6ffef85ffe5f5;
assign w_fix[46]='hfffe330012cd00190bfffd07ffeef3;
assign w_fix[47]='hfff2d7000e7b001887000771fff71c;
assign w_fix[48]='hfff8ad000952000b2fffff9bfff84e;
assign w_fix[49]='h0001c0001512000375fff088ffecb3;
assign w_fix[50]='hfffeff000ed4fff69bfffc1cfff0da;
assign w_fix[51]='hfff73500016dfff9a80007ec000111;
assign w_fix[52]='hfffff9ffff4c000027000352000009;
assign w_fix[53]='hffffebfffa1cfff8fafffc6100002e;
assign w_fix[54]='h000030000642fffe57fff3d1fffdb1;
assign w_fix[55]='hffff7bfffd88fff5b80007fcfffcf4;
assign w_fix[56]='hfffe2ffff9e2000a99ffe47effff73;
assign w_fix[57]='hffffcf000d9efff6fb0005d3fffd86;
assign w_fix[58]='hfffcbb00134bfff77d001751000059;
assign w_fix[59]='hffff04000e1e000187fff1fffffda7;
assign w_fix[60]='hfffd43000debfffb63fff0dafffe76;
assign w_fix[61]='hfffcbb000e15fff44effe809fffe9c;
assign w_fix[62]='hfffe36fffbc30016b7ffecfafffef8;
assign w_fix[63]='hffff49ffe7d40000080009a7fffe94;
assign w_fix[64]='hffff8c00021900041c0012d1fffe20;
assign w_fix[65]='hffff5200037d000953001368ffff0d;
assign w_fix[66]='hffff5d00006600031c001806ffffb3;
assign w_fix[67]='hfffe2cfffeff00015d0009b9fffef7;
assign w_fix[68]='hfffc73fffff00005b7fffe95fffe3c;
assign w_fix[69]='hfffd290014150012b300088efffd64;
assign w_fix[70]='hfffbfe001e85ffef1d000ffafffc75;
assign w_fix[71]='hfffe4e001fee0003fa0003edffff34;
assign w_fix[72]='hfffe1c000673001b05ffeffefffccf;
assign w_fix[73]='hfffdbb000a2300070bfff7eafffd8d;
assign w_fix[74]='hfffd06001087000515fffdcefffeaa;
assign w_fix[75]='hfffc840004e0fffbf9ffe97dfffeea;
assign w_fix[76]='hfffd87fff6a7ffff55ffe4b2fffe4a;
assign w_fix[77]='hffff4a000207fff92cfffbaeffffdc;
assign w_fix[78]='hffff71fffa86fffed400016e0001f3;
assign w_fix[79]='hfffa94fff1dbfff5fc000762fffd37;
assign w_fix[80]='hfff649ffe35afffb850006c7ffe46e;
assign w_fix[81]='h000381ffe79afff3d400036cfffd10;
assign w_fix[82]='hfff2c4ffe555fff5b4001a15ffd642;
assign w_fix[83]='hffea28fff55bfff105001893ffef7d;
assign w_fix[84]='hffef85000b4affebfa000a97fff192;
assign w_fix[85]='hfff512000064ffed63000e4cfff6e4;
assign w_fix[86]='hffeb32fff499ffef9e000e82fff64e;
assign w_fix[87]='hffed9f0009c7fff67b00044ffff251;
assign w_fix[88]='hfff97400005cfffe320006c7ffe47a;
assign w_fix[89]='hfff8e4fff108fffacc0004c9fff1e0;
assign w_fix[90]='hffff84fff79ffffb87fffebb000882;
assign w_fix[91]='hfff963ffede8fffbb300044b000b65;
assign w_fix[92]='hfffb9bfff760fffaa5000287000d38;
assign w_fix[93]='hfff3e6ffe94afff57d00057efff041;
assign w_fix[94]='hfff22a0002a1fff2a3000de6fff00c;
assign w_fix[95]='hffed55fffafeffefd9001889fff183;
assign w_fix[96]='hffe77afffb1fffee0f0008aafff796;
assign w_fix[97]='hfff16efff21dfff352000ec6ffe4b1;
assign w_fix[98]='hfff5bafff193fff3b6000d41fffb73;
assign w_fix[99]='hfffd83ffeb89fff67c000682000459;
assign w_fix[100]='hfffeb5ffe042fff9d50006e9fffbfd;
assign w_fix[101]='hfff6c1ffcf8ffffce8000878ffe36e;
assign w_fix[102]='hfffd11ffe179fff6d3000ba2ffec17;
assign w_fix[103]='h0004fffffae7fffe5700005200083f;
assign w_fix[104]='hffff45fffcf9000bcbffff9affff62;
assign w_fix[105]='hfffd2ffff292001eed001503000bed;
assign w_fix[106]='h00017dfff28e003cec0008fdffffa8;
assign w_fix[107]='h0011f3ffe983001c570005910008ff;
assign w_fix[108]='h0012780018df000100000620001051;
assign w_fix[109]='hffe98f000ca3fffd430003f80004c7;
assign w_fix[110]='h00054dfffc7dffe5d6ffe45e001216;
assign w_fix[111]='h001c02ffe9f4ffef6efff285002ce0;
assign w_fix[112]='h000135fff67afff270ffefb8002cce;
assign w_fix[113]='hfff1e3fff82e00025cffe289001d34;
assign w_fix[114]='h0010ba002b4effd676ffe2dd001526;
assign w_fix[115]='h000b03fff6c6ffdbc6fffe39000ecd;
assign w_fix[116]='hfffdfbfffebb000147ffff300005c0;
assign w_fix[117]='hffe60900082efffdc2001b8efff33e;
assign w_fix[118]='hfff8d9fff9b800078c000df7fff327;
assign w_fix[119]='hfff4feffef5f00073100078800033f;
assign w_fix[120]='hffd8d1ffe806001767000c70001760;
assign w_fix[121]='hffe7c1ffefc1fff753001e26fff4f2;
assign w_fix[122]='h0001c8ffe92a00162dfffce9fff5db;
assign w_fix[123]='h000d7b000035001d3d0001a7ffebfc;
assign w_fix[124]='hfff9f6001a26fffeaefff9f5ffe95b;
assign w_fix[125]='h0001af0013b5fffba4fffe66ffebec;
assign w_fix[126]='h000abc001076001580000ef7ffebda;
assign w_fix[127]='h000d62000571000878001ac0ffffb5;
assign w_fix[128]='h000ffaffea93000928000fe60011f0;
assign w_fix[129]='h00096ffff3a00001ad000366000d3a;
assign w_fix[130]='h00001afffd7ffffe07fffdcc000071;
assign w_fix[131]='h000078fff98f00046bfff4ecfffda2;
assign w_fix[132]='hfffe3efffac400030ffff3f7fffeae;
assign w_fix[133]='hfffdfaffe955000811fff11dfffcae;
assign w_fix[134]='hfffd1300179afff29c001470fffc07;
assign w_fix[135]='hfffb16000a950006de0017fafff912;
assign w_fix[136]='hfffd08ffe8240009f2000f28ffff34;
assign w_fix[137]='hfffc75ffe30e000559fff3dcfffd69;
assign w_fix[138]='hfff946ffebd3000fc5ffee6efffd9c;
assign w_fix[139]='hfff9b7fff406000a26ffed2afffdc0;
assign w_fix[140]='hfff89f000cf3fffa22fff9ae0001a7;
assign w_fix[141]='hffffa6ffec56fff42dfff93afffe16;
assign w_fix[142]='hfffeeefff8c9fff878fff6d7ffff41;
assign w_fix[143]='h0000b40002f1fff43c000121fffece;
assign w_fix[144]='h000062fffb2bfff0e3fffc40fffeee;
assign w_fix[145]='hffff20fffb80fff018fffe42fffbc5;
assign w_fix[146]='hffff7dfff886fffce3000254fffc29;
assign w_fix[147]='h000565ffec7a00045900136afffd8c;
assign w_fix[148]='hfff665fff55c0015af000865fffbe1;
assign w_fix[149]='hfffbb1000b8f00152a0008540003a9;
assign w_fix[150]='hfffa970011920003eb00070500020d;
assign w_fix[151]='hfffb6d000028000bc6fff7dffffef4;
assign w_fix[152]='hfffe390003b5000516fff5360000cb;
assign w_fix[153]='h0000100004ecfffb5b000e90fffd7b;
assign w_fix[154]='hfffe65fff5040000ae000ec0fffd75;
assign w_fix[155]='hfffee3fffc4a000842fffaf3fffdca;

endmodule