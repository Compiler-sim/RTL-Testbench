module wf_buffer #(
  parameter D_WL = 24,
  parameter UNITS_NUM = 5
)(
   input [7:0] addr,
   output [UNITS_NUM*D_WL-1:0] w_o
);


wire [D_WL*UNITS_NUM-1:0] w_fix [0:155];
assign w_o = w_fix[addr];
assign w_fix[0]='h000015000144fffe7effffe6001261;
assign w_fix[1]='hfffee70009b1fff46cfff9390021e5;
assign w_fix[2]='hfffb94fffa47000086fff85b000d63;
assign w_fix[3]='hfffd85001133ffe9eefff667fff89a;
assign w_fix[4]='hfffe2c0009b6fffe07fffbd8ffece6;
assign w_fix[5]='hfff9fe001e86fffeeffffb5afffe00;
assign w_fix[6]='hfff90c0027e0000d97000097000bd0;
assign w_fix[7]='hfffe90001d30000c06fffb31001c60;
assign w_fix[8]='hfffd830020c400029bfff84b0006fa;
assign w_fix[9]='h0000c5000de5fff6c1fff753fffda9;
assign w_fix[10]='h0001580009e50009630001a3ffe5fc;
assign w_fix[11]='hfffef3000451000e9a00005f000229;
assign w_fix[12]='hffff9bfffea2fff743fffff6fffe9b;
assign w_fix[13]='hfffcccfffe78fff984ffff34fff5de;
assign w_fix[14]='hfffe67ffff10fffecdfffd26fff98b;
assign w_fix[15]='h00004affec6a00092ffff678ffff43;
assign w_fix[16]='h00011cfff12b0010fbfff403fffac1;
assign w_fix[17]='hfffc6f0005ab0005d8fffc49fffef2;
assign w_fix[18]='hfff796fff18afff57afff587fff0fc;
assign w_fix[19]='hfffc08ffea390008f7fffa15000072;
assign w_fix[20]='hfffe95fff671fffd52fffd0200028a;
assign w_fix[21]='hfffbf8000d2dfff194fffe50000159;
assign w_fix[22]='hfffa3c000cc4000541fffed6fff873;
assign w_fix[23]='hfff8c2ffefc5fffc38ffffc7fffa86;
assign w_fix[24]='hfffc6effff57fff3bffffeb40007fe;
assign w_fix[25]='hfffe5dfffc7dfffff9fffe9dfff7c8;
assign w_fix[26]='hffff0f000483ffffdd0001f50001b4;
assign w_fix[27]='hfffdb20018c0fffa88000fda001305;
assign w_fix[28]='h00076effec04ffef37002aa4001b51;
assign w_fix[29]='hffea4dffe814ffeab8002deb001ce3;
assign w_fix[30]='h001a58fff735fffc250032f90014ac;
assign w_fix[31]='hfff397fffe31fffb94003afa001399;
assign w_fix[32]='hffef2b000d2700044f000d4f000b2e;
assign w_fix[33]='hfff35c00143200034f00051e000489;
assign w_fix[34]='hfff0ca00136ffffbc0fff5660006d2;
assign w_fix[35]='hffed4400034ffff87500062e0005ba;
assign w_fix[36]='h000390001db900050effedbb000120;
assign w_fix[37]='hfffdfe0022cf000602ffdd93000149;
assign w_fix[38]='hfffd820016140005f8fff66c000456;
assign w_fix[39]='h00003d00131500085bfff950ffffa1;
assign w_fix[40]='hfffb9a000b1d000502fffba4000129;
assign w_fix[41]='h00072700113c0006cafffb470000d6;
assign w_fix[42]='h00121b000d7500022e0008030003fe;
assign w_fix[43]='h0006560013180006330019b8000776;
assign w_fix[44]='hffee01fff8460000b2000da800034c;
assign w_fix[45]='hfff6be00012000017b000a380003cf;
assign w_fix[46]='hfffce50007c4000979000bf8000b29;
assign w_fix[47]='hfff8d2fffc7d0006bbfff9cb00098d;
assign w_fix[48]='h0003cdfff1c1fffeeffffbe600063a;
assign w_fix[49]='h000db6000f5dfff4e00000cd0003fb;
assign w_fix[50]='h00082b0011dffff253fff994000988;
assign w_fix[51]='hfffab5fff65cfff9c5fffabf0005f0;
assign w_fix[52]='h0000030001f8000006000a9afffff9;
assign w_fix[53]='hffffd9000534fffb52003034000034;
assign w_fix[54]='hffffabfff11c00090400088dfffe31;
assign w_fix[55]='hffff98ffe6e1fff5c0002673fffdf6;
assign w_fix[56]='hffff44fffcc4000b6b000825ffff20;
assign w_fix[57]='hfffeeefff94000003f00274bfffe66;
assign w_fix[58]='hfffd10000a12fff1d1000e6dfffef3;
assign w_fix[59]='hfffe880010ddfff566000a22fffddc;
assign w_fix[60]='hfffda2000b87fff39afffb5afffe40;
assign w_fix[61]='hfffe36fff642fff6e2000852ffff17;
assign w_fix[62]='hffff40ffe7af000171000193ffffb2;
assign w_fix[63]='hffff8fffee6afff71d000556ffff66;
assign w_fix[64]='hffffbbfff5f6ffff3f0013a2ffff00;
assign w_fix[65]='hffffb0fff95900045d00186fffff63;
assign w_fix[66]='hffffcbfff853fffe55001bc3ffffe8;
assign w_fix[67]='hffff52fff51cffff8bfffe2dffff9e;
assign w_fix[68]='hfffdc400042d00021ffff276fffef0;
assign w_fix[69]='hfffe1b0004550001e900023bfffe83;
assign w_fix[70]='hfffd0a000030ffe870000612fffd55;
assign w_fix[71]='hfffe1ffffe0efff6a900070fffff0a;
assign w_fix[72]='hffff34000490fffeee00021cfffe77;
assign w_fix[73]='hffff16fffd7dfffb8d000152fffecf;
assign w_fix[74]='hfffecdfff854ffff23000bc8ffff9e;
assign w_fix[75]='hfffe9ffff903fffdc7000fe0ffffef;
assign w_fix[76]='hfffec3fff97ffffcda00126dffff6c;
assign w_fix[77]='hffffc7fff5c9fffce6000e1e000013;
assign w_fix[78]='h0001570006d300003dfff80a0000b8;
assign w_fix[79]='h00068c0013f3fff7e2fffe14001235;
assign w_fix[80]='h00089d001003fff73affcdd9001ee2;
assign w_fix[81]='h0015e4001086ffeaebffe7840021cc;
assign w_fix[82]='h000f9b000d56fff65d0027f2002115;
assign w_fix[83]='h000968000e380016b1001f36001dd1;
assign w_fix[84]='h000cbe001ad9000777002a2e000e45;
assign w_fix[85]='h000d5a001085000a2a002234000986;
assign w_fix[86]='h0003010010d6fff8d400203e000543;
assign w_fix[87]='h000e8a000b70ffff8f00117f000588;
assign w_fix[88]='h000f12fff795fffd2f002328fffcf1;
assign w_fix[89]='h00084f0001b8000333001786fffb52;
assign w_fix[90]='h0007ca000783fffc7c0009e5000140;
assign w_fix[91]='h000450000aedfff92f0010d300004e;
assign w_fix[92]='h0005b6000935fffbebfffb24000304;
assign w_fix[93]='h00042d000ec8fffa17ffed21fffeb5;
assign w_fix[94]='h0004c5001c4dfffb9100065d000310;
assign w_fix[95]='hfffe5d001af5000668000e3d00093e;
assign w_fix[96]='h000542000b87ffeea0fff3290004a6;
assign w_fix[97]='h00136300075bfffe4cffe99d00037f;
assign w_fix[98]='h0002ba0001cdfffae0000b7a001259;
assign w_fix[99]='h000218fffceefff540000c42001507;
assign w_fix[100]='h0001f400009c000054fff51d000c0e;
assign w_fix[101]='h0005240003510002960003650008d2;
assign w_fix[102]='h0004b4000364fffddd0006f30015b7;
assign w_fix[103]='h0001fd0000e0ffff58000156001479;
assign w_fix[104]='h000381fffa530010320003c600110a;
assign w_fix[105]='h000024fff22600291b0010ac001dc1;
assign w_fix[106]='h000df7fff136002ae100119a0005fc;
assign w_fix[107]='h001774ffdb8c003f4d000c3f000675;
assign w_fix[108]='h000fa2001edd003a11000a310017f4;
assign w_fix[109]='hffef7c0008ab0026d800136e000ed9;
assign w_fix[110]='hfffb3fffecb500233a00043a000b61;
assign w_fix[111]='h0014bcffe19cffed70000abd002bb0;
assign w_fix[112]='hffead4ffede2ffeba8000029001ca7;
assign w_fix[113]='hffd63a0005b0fff9d0fff85e001e54;
assign w_fix[114]='hfff67000282bfff8e900042b000409;
assign w_fix[115]='h001f40fff352fff3e800071e0005e7;
assign w_fix[116]='h001057fff3b400078d0000ed000d01;
assign w_fix[117]='hffffbd00007500040f0004db001083;
assign w_fix[118]='h00024efff4db0013cc00099400068c;
assign w_fix[119]='h000026fff3e6000510000b390013dc;
assign w_fix[120]='hfffb20fff61d000f20000c980016d1;
assign w_fix[121]='hfffccdffffc000194b000d6b000019;
assign w_fix[122]='hfff3d5fff44f00147f0010080002a5;
assign w_fix[123]='hfff46afffd51ffef3b000fdf000752;
assign w_fix[124]='hfff36c0000b60001b10005e0fffec1;
assign w_fix[125]='h000104fff834000cb100038dfffeb7;
assign w_fix[126]='h0012ff000c6c0005c700047afffc8c;
assign w_fix[127]='hfffdda001050fff7ed000b070006b0;
assign w_fix[128]='h0004e0000422fff9810009ec00148f;
assign w_fix[129]='h0000820000ea001cd7ffff2a000ce1;
assign w_fix[130]='h00001bfffc79ffff59fffe4d000090;
assign w_fix[131]='h000069fff56e001eb6000245fff736;
assign w_fix[132]='hffffdaffed27fff2e8fff380fff055;
assign w_fix[133]='hffffd1ffdafdffdfe4fff384fff124;
assign w_fix[134]='hfffec600191efff182000947fff8c8;
assign w_fix[135]='hfffd700003bcffe7e3fff931fff76e;
assign w_fix[136]='hfffec8ffeacbffff60000badfffe06;
assign w_fix[137]='hfffd79ffe589001462000a67fff788;
assign w_fix[138]='hfffc3ffff5ca000a08fff866fffc40;
assign w_fix[139]='hfffe95fffb4d0014f4ffeb5ffffb20;
assign w_fix[140]='hffff9c00155c0000230000ecffffdb;
assign w_fix[141]='h00006dffeff5ffd9a8000355fffd8d;
assign w_fix[142]='h000000fff675ffea4f000048fffef1;
assign w_fix[143]='h000054ffff30ffe84c000295fffc6f;
assign w_fix[144]='h00004efff83effe9e0fffda7fffc8a;
assign w_fix[145]='h000072fff531fff5f50003cefff5a5;
assign w_fix[146]='h00004dfff5940015e40006adfff23f;
assign w_fix[147]='h00019affebe900204e0012a7fff6bd;
assign w_fix[148]='hfffcacffec67001448fff98afff5ab;
assign w_fix[149]='hfffdd1fff9dd00154efffb39fffb8f;
assign w_fix[150]='hfffea0ffffd9fff6c0fffa82fffc64;
assign w_fix[151]='hffff7cfffe75ffe790fff882fffb1b;
assign w_fix[152]='hffff810005d1fff79bfff7cdfffd91;
assign w_fix[153]='hffffdb00086afffe75000ceefff9ea;
assign w_fix[154]='hffff62000469fffb9d001681fff868;
assign w_fix[155]='hfffffd000358fff9c4fffc95fff875;

endmodule