module wg_buffer #(
  parameter D_WL = 24,
  parameter UNITS_NUM = 5
)(
   input [7:0] addr,
   output [UNITS_NUM*D_WL-1:0] w_o
);
//156*5=26*30
wire [D_WL*UNITS_NUM-1:0] w_fix [0:155];
assign w_o = w_fix[addr];
assign w_fix[0]='h0002b900109ffff8440004790003ee;
assign w_fix[1]='hfffe7400167bfff888000a700035a3;
assign w_fix[2]='hfff822fff927001678002b42003302;
assign w_fix[3]='hffeff70013f4ffe96f001249002257;
assign w_fix[4]='hfff3400009abfffb050016fa001277;
assign w_fix[5]='hfff0ba002131000412000fa3fff935;
assign w_fix[6]='h00064f001d360019d20016eaffe841;
assign w_fix[7]='h000b280014f70017540015f9fffd81;
assign w_fix[8]='h001405000d40001233001a3100156f;
assign w_fix[9]='h00167a000424000f69001593000f5c;
assign w_fix[10]='h0010120000a000176e0015dbfffa05;
assign w_fix[11]='h000c2e000c79000a2b0012fbffd96d;
assign w_fix[12]='h000db100025bfff408000624fffc49;
assign w_fix[13]='h000e780005880000a1fffccbfff031;
assign w_fix[14]='h0015f900042b000933fffa06ffe496;
assign w_fix[15]='h001b2afff17a0005a3ffeb2efff566;
assign w_fix[16]='h001b61ffeb1e0016a6ffe74200010a;
assign w_fix[17]='h00163c000f04002a21fffcd5ffec08;
assign w_fix[18]='h001156fff6040018c4fffec7fff906;
assign w_fix[19]='h0024dffff4d60016430006050000a1;
assign w_fix[20]='h0029cf000aceffecb70004fffff55d;
assign w_fix[21]='h00202e001234ffd8b7000463fffdb9;
assign w_fix[22]='h002314000ad0ffcefa0009cefff8d6;
assign w_fix[23]='h0027110008eaffd29e000ebafffad2;
assign w_fix[24]='h00265c000fbeffc8f3000cad0005ab;
assign w_fix[25]='h001528001435ffb8bbfffe46fff887;
assign w_fix[26]='hfffa5efffd3d00001d0006a8000117;
assign w_fix[27]='h00071cffcdc9fff502000cd20009a9;
assign w_fix[28]='h00049dffd835fff624fffdf6000d6d;
assign w_fix[29]='hfffd80fff29bfffd750017d9000e5e;
assign w_fix[30]='h0031cdffd60fffee840029c5000aff;
assign w_fix[31]='hfffe3e00090bfff2b20024ab00090f;
assign w_fix[32]='hfff5fd00023efff1ec000ec900069a;
assign w_fix[33]='h0005d60004effff5f3000bd800064c;
assign w_fix[34]='hfff80efff321fffd750005ba000704;
assign w_fix[35]='hfff0f5ffd34affef35000094000694;
assign w_fix[36]='h00061fffe200ffd916fff69c000355;
assign w_fix[37]='hfff28bffe84fffea4dfffacc000584;
assign w_fix[38]='hfffbe8ffeff40002a7fffe3200042b;
assign w_fix[39]='hfff8de0005f60010dfffff0b0000f1;
assign w_fix[40]='hfff631000f9f000dc5000786000788;
assign w_fix[41]='h00135ffffe83ffff4e00100b000eb5;
assign w_fix[42]='h0019670013e0ffefbe0013fc001173;
assign w_fix[43]='h000319000d07ffee6600080e00110e;
assign w_fix[44]='hfff2f20004cd0006b8000c0400194e;
assign w_fix[45]='h000114ffdd7400037a00105d001a63;
assign w_fix[46]='h0000c7fff60b000f780014f3001966;
assign w_fix[47]='hffed5dffec56001a040014ce001bfb;
assign w_fix[48]='hffedbffff288001b1a001aa3001dcd;
assign w_fix[49]='h000cd1ffe92300041900174f0021c4;
assign w_fix[50]='h000887ffeda1000272001e1900254e;
assign w_fix[51]='hffe52c0010c1000ed8002273002a6a;
assign w_fix[52]='hfffea500013afffec4000145ffff3d;
assign w_fix[53]='hffffffffdba20003b5000af3fffe00;
assign w_fix[54]='h000c4dffdd2b0012d5fff813ffff02;
assign w_fix[55]='h000510ffe256001357fff04ffff7a6;
assign w_fix[56]='h000abbffd4120020b0ffedee0003b6;
assign w_fix[57]='h000ea6ffd57a000c7600016cfff8bf;
assign w_fix[58]='h000c77ffe98a0009a0001881fffbbc;
assign w_fix[59]='h0001fbfff23600082f000228fffddc;
assign w_fix[60]='hfffaf9fff6d8000712000ea1000195;
assign w_fix[61]='hfff684ffe93c0019bd001f3e000c31;
assign w_fix[62]='hffff55ffefbe001bb700196b00107a;
assign w_fix[63]='hfffac000008f000dda000a47fffd53;
assign w_fix[64]='hfff961fffd1b0008c0000e90fffe4c;
assign w_fix[65]='hffff090010bafff7720003acfffa43;
assign w_fix[66]='hfff508001769fffb6cfffee1fffc5f;
assign w_fix[67]='hffefc8fffbfb000a36000548fff9aa;
assign w_fix[68]='hffef94ffeed8001272001276fff93d;
assign w_fix[69]='hffffe700035d000dc1fffdc2fff7a6;
assign w_fix[70]='hfff8ed0003abffffc7ffe823fff753;
assign w_fix[71]='hfff3a80008e40017ddfff1c9000038;
assign w_fix[72]='hffeb2d000c35000d34000425000413;
assign w_fix[73]='hffec890015cdfff342000f41fffa6c;
assign w_fix[74]='hffec580016f2ffe9b90011bdfffc50;
assign w_fix[75]='hfff3b900054ffff28bfffad70001a3;
assign w_fix[76]='hffee39fffba5fff7a000219900023a;
assign w_fix[77]='hfff04dfff924ffea840026a4fffae7;
assign w_fix[78]='hfff8ad000449fff50bfffea7fff76a;
assign w_fix[79]='hffec82000997fff41e000720fff38d;
assign w_fix[80]='hffd4e9fff53effffe4000e7bffe3c9;
assign w_fix[81]='hffcfaa00001cffdcdbfffffcffe93f;
assign w_fix[82]='hfff5bbfff66b001404001dbdffe92e;
assign w_fix[83]='hfff7e1fff54a00076fffef67ffe900;
assign w_fix[84]='h0010a3000be40011540016bcfff911;
assign w_fix[85]='h000d980026a2000e36000d26002adb;
assign w_fix[86]='hfffbf30009a3fff58c001ca00018ca;
assign w_fix[87]='hfff3df000239fff3d70023aa000122;
assign w_fix[88]='hfff11900065efffa87001b26fff44b;
assign w_fix[89]='hfffe82001460ffea14000f460004a3;
assign w_fix[90]='hfff27d000635ffe221000964fffbc8;
assign w_fix[91]='hfff550000d8cffe4ddfffcb6ffff15;
assign w_fix[92]='hfff31b000fbcffe4a2fff5f4fff591;
assign w_fix[93]='hfffc46000f82ffff22001410ffec62;
assign w_fix[94]='hfffa1b000f0c00077d000d78fff171;
assign w_fix[95]='h0012ce000552001560000d82fff547;
assign w_fix[96]='hffeebc0012bc000bd4fff88fffeddc;
assign w_fix[97]='h0002010016500009a20021a90002a3;
assign w_fix[98]='hffff63fff4d2fff1500016eeffe90f;
assign w_fix[99]='hffed7fffe7d3ffcf5c000a83ffd1d2;
assign w_fix[100]='hfff23bfff3feffcd96fffdd1ffd0dc;
assign w_fix[101]='h001406fff3f3ffda73000976ffcd18;
assign w_fix[102]='h000e6fffe19dffe17f000ab0ffc55c;
assign w_fix[103]='hffe320ffe14affd0840002b8ffba3c;
assign w_fix[104]='h00096efff90fffed8d000055000487;
assign w_fix[105]='h000902000684ffe7f6000890002b9b;
assign w_fix[106]='h002e9d001cfeffd888001a86003bbf;
assign w_fix[107]='h002b4b001925ffe6ca000c0b003bfa;
assign w_fix[108]='h00008400456800008700019a001bb6;
assign w_fix[109]='hfffedc002e1bfff84efffe9b001936;
assign w_fix[110]='hffe08f00067b001e37000516fff18c;
assign w_fix[111]='hffe15e00036c00129d0003f0ffd025;
assign w_fix[112]='hffee8e000e87000c0afffd93ffde7f;
assign w_fix[113]='hffffec001f11001d7500031dfff8ab;
assign w_fix[114]='h000976002c640032ff000d280014e7;
assign w_fix[115]='hfff57bfff72200127a000531ffeeb9;
assign w_fix[116]='h000dabfffaf40013230004c00001be;
assign w_fix[117]='h000736ffefe0fff86d000b90fff247;
assign w_fix[118]='h0000d4ffe963fff6680005dffff33d;
assign w_fix[119]='hffe3ccfffa81fff43efffb96ffff04;
assign w_fix[120]='hfff194fff4ec0009770000c0fff975;
assign w_fix[121]='hffeae8ffe901000b80001133ffff10;
assign w_fix[122]='h00170cffed99ffe2df000913000f3f;
assign w_fix[123]='hfffe90fffbf4ffee290004d8000902;
assign w_fix[124]='h000d82ffff290019aafffc7500082d;
assign w_fix[125]='h001b82ffeff600087b00079800018d;
assign w_fix[126]='h0000f3fff2baffff9e0009b9fffc67;
assign w_fix[127]='hffd3affffd79ffdeef000bbcfffa96;
assign w_fix[128]='hffe844fffda20006b0000a39000311;
assign w_fix[129]='h002c96ffeabd0022920004880012f6;
assign w_fix[130]='h000018fff958fffff6000274ffed6b;
assign w_fix[131]='hfffd42fff95afff1a4002a06fff394;
assign w_fix[132]='hfff7ff0013bcffdbd400243bffee8e;
assign w_fix[133]='hfffbe7000dd2ffe1a6001233fffd55;
assign w_fix[134]='h000463003d42ffcc3c00363effef58;
assign w_fix[135]='h00060a00307fffda7cfff6cafff497;
assign w_fix[136]='hfffe7d0017ceffedcafffd70ffe29d;
assign w_fix[137]='h00011200071c0002f1fff9a2ffe461;
assign w_fix[138]='h0003330007c4fff911fffd50ffd388;
assign w_fix[139]='hfffd34001562fff76300160fffdc37;
assign w_fix[140]='hfffb450016730001d0000c80ffd997;
assign w_fix[141]='hfffdddfff234001438fff915ffdb9f;
assign w_fix[142]='hfffedcfffaf8ffffc80001b6ffe6fc;
assign w_fix[143]='hffff58fff0f50007e4fff3ccffe1fd;
assign w_fix[144]='hfffe65ffe269000cdbfff6f9ffde33;
assign w_fix[145]='hffff30ffeea1000782000aa4ffee7a;
assign w_fix[146]='hfffd96ffe627fff9b8000777fffa6a;
assign w_fix[147]='hfffc20ffec48fffa5f0011b4ffeafb;
assign w_fix[148]='hfffcf5fff7ac00135f0002abfff3e2;
assign w_fix[149]='hfff70d0005d9001fdf001208ffe5f2;
assign w_fix[150]='hfffae800145e000a63000a20ffd854;
assign w_fix[151]='hfffe8efffe210000a3000385ffd93b;
assign w_fix[152]='hfffdc9fff450000265fffd7dffd1b6;
assign w_fix[153]='hfffa9a0000780007490018c9ffcc55;
assign w_fix[154]='hfffac0ffff92ffe6e1001c7fffd141;
assign w_fix[155]='hfffee5ffedaeffe174fff8e9ffec00;

endmodule