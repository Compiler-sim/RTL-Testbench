module ri_buffer #(
  parameter D_WL = 24,
  parameter UNITS_NUM = 5
)(
   input [7:0] addr,
   output [UNITS_NUM*D_WL-1:0] w_o
);

wire [D_WL*UNITS_NUM-1:0] w_fix [0:179];
assign w_o = w_fix[addr];
assign w_fix[0]='h0001ac000e83001948ffe36bfff8d5;
assign w_fix[1]='h00021500235200023afff1ce001ff7;
assign w_fix[2]='h000a85ffeea90004f0fffbd5fff9cd;
assign w_fix[3]='hfff2aefffc060025fe0008c800075a;
assign w_fix[4]='hfffdb3000a5e000653ffeea00030b1;
assign w_fix[5]='h0009ddfffc34fffa3dfffe79ffe33a;
assign w_fix[6]='hfff2480000ea00047dfffbb1ffe85d;
assign w_fix[7]='hfffe6d00154affecfc0003e5fffd26;
assign w_fix[8]='h00108b002bc3001464000280fff8ff;
assign w_fix[9]='hfffe2700006a00139c0000fe00003f;
assign w_fix[10]='h0001380008ac000743fffbdd000920;
assign w_fix[11]='h000140ffdc6c000081ffe20e000c77;
assign w_fix[12]='hfffaf90008d80018a7fff924fffb1a;
assign w_fix[13]='h001023000a20ffe9b9000a6900124d;
assign w_fix[14]='h0002a0fffd9e00017e000008ffff39;
assign w_fix[15]='hfffbdd000b320000cb0004d50020cb;
assign w_fix[16]='hffe9ad00067c0011e0fffa75ffeb32;
assign w_fix[17]='h00065a000b2cfff14bfff9b8000e0c;
assign w_fix[18]='h0007eb0010ee00008a0002990009c7;
assign w_fix[19]='h0000a1fff6c0000021000226002659;
assign w_fix[20]='hfffabfffeeaffffb9efff8e6ffe154;
assign w_fix[21]='hfff6bcffe8e5fff634fff76effe7b1;
assign w_fix[22]='hfff0c700034b000155fff8f4ffee88;
assign w_fix[23]='hfffbd800077f000cd7fff719fffdec;
assign w_fix[24]='hfff9550005b0fff470fff437ffda8a;
assign w_fix[25]='hfffd9effd9d1fffcbc001662ffc5f2;
assign w_fix[26]='hfff794fff44e0007b3fffcf7000ec7;
assign w_fix[27]='h00021e0008e5fffbe20014cd00213d;
assign w_fix[28]='hfff8950002f4000d17fffd41ffff1d;
assign w_fix[29]='h000143fffdac0000ea000570000401;
assign w_fix[30]='h000fa0fff509fff941fff150000f7b;
assign w_fix[31]='hfff355fff886fffbf60023a7fffe6a;
assign w_fix[32]='h00093dffffdafffb34001049000d5b;
assign w_fix[33]='hfff36f0000a9000871ffe8cb0013ab;
assign w_fix[34]='h00009efff83ffffef3000dcffffbae;
assign w_fix[35]='hfff7c2000144fffe9affe3e6fff815;
assign w_fix[36]='h0001d400130f0002660003120000f3;
assign w_fix[37]='h000042000f59000250fff7a1fffd5a;
assign w_fix[38]='hfff7fb0003100009e6fffe92fff7b5;
assign w_fix[39]='hfffdc2ffea02fffd1d00189b000ad7;
assign w_fix[40]='h000039fff202fffd1c000ab100031f;
assign w_fix[41]='h000f900016770003c3ffe545000b07;
assign w_fix[42]='h00074bfff00b00015200136b000875;
assign w_fix[43]='hfffc2b0006b0fffeb700002affeb1e;
assign w_fix[44]='hfffeaffffe31fffefe000e94000250;
assign w_fix[45]='h000c6dfffa180002990021510003b9;
assign w_fix[46]='h001defffec9900023e000672ffff66;
assign w_fix[47]='h0000fffff7e2fffaf800154afffcc0;
assign w_fix[48]='h0009e0fff50ffffcdd001098000083;
assign w_fix[49]='h000631fff91dfffd17001823fff69a;
assign w_fix[50]='hfffdc9fff37bfffe210003120014d8;
assign w_fix[51]='h000a45fff2ddfffad6fffbec0006b5;
assign w_fix[52]='h0000c900200e00084d00168c00232a;
assign w_fix[53]='hffffb5fff41ffffcd20033000007bc;
assign w_fix[54]='hfff9f4ffede9000154fff836001694;
assign w_fix[55]='h00037effff37fffd77ffda66ffffd7;
assign w_fix[56]='h000d1effff2f0001f0000d990002ed;
assign w_fix[57]='hfff7fb000ce80004900008edfff137;
assign w_fix[58]='hfffec9ffec11fffd620032ae0008f7;
assign w_fix[59]='hffffec00065300013a000606000069;
assign w_fix[60]='hfffc1a000d03fff1e2ffdb600000d6;
assign w_fix[61]='hfffec8000771fffd980012a00001ad;
assign w_fix[62]='hffffa3ffe354fff9a1ffff2c000207;
assign w_fix[63]='h00012000052a0002ceffd84ffffa08;
assign w_fix[64]='hffff7e000a9e000478000cb3fffffc;
assign w_fix[65]='hfffc79fffe64fffa5cffd2bbfffe32;
assign w_fix[66]='h0000b2000e2fffeec3ffe1e6fffcfe;
assign w_fix[67]='h00009e00016b00056ffff5d30000c0;
assign w_fix[68]='h000a310014f500072f0009930000ff;
assign w_fix[69]='hffff99fff056000836fff960fffea5;
assign w_fix[70]='hffffb200014600000d000010000198;
assign w_fix[71]='hffff88fffb76000002ffff46fffff0;
assign w_fix[72]='hffff3ffffb2900062bffef87ffffec;
assign w_fix[73]='h0000d3fffca70015550003460004cf;
assign w_fix[74]='hffffa7ffff8cfffe51000440fffff9;
assign w_fix[75]='h000438000366000eb30027a80008f8;
assign w_fix[76]='hfff8ecffff230012f2ffe95dfffd08;
assign w_fix[77]='h0000bc000af5fff6aefff5dfffff5c;
assign w_fix[78]='hffffb6ffec69000941fff8ad0001c3;
assign w_fix[79]='h0000710006090002bd000daa0001e0;
assign w_fix[80]='hfffd090009c9fff1b30004030002ca;
assign w_fix[81]='hfffa8dffe45c000543ffe5f9fffc0d;
assign w_fix[82]='hfffeec001678fff315ffe48a000220;
assign w_fix[83]='h0001c9000a99fffd54000751000141;
assign w_fix[84]='h000133fff953fff8c80000bdffff26;
assign w_fix[85]='hfffe87ffed4bfffb1cffe56efffea2;
assign w_fix[86]='hfffe5afffc1b000a2cfff908ffff56;
assign w_fix[87]='h0002560004800008a0fff859ffff47;
assign w_fix[88]='h000063000392fffe04ffff8affffa1;
assign w_fix[89]='h00011900066dfffea800055100006b;
assign w_fix[90]='h0010ee000e92fff755ffcd17000d2c;
assign w_fix[91]='hfffd4b00079f0017e8fffe1f00195d;
assign w_fix[92]='hfff9fd000adb000bf2000e2b0015de;
assign w_fix[93]='h0003cafffda3fffff50008e4000e3b;
assign w_fix[94]='h000151000df6000ffa00013e001099;
assign w_fix[95]='h0002b1fff025ffee39000435ffe854;
assign w_fix[96]='h00073cffefd1fff24affe8cc0006bd;
assign w_fix[97]='h000033ffed7bfff9d0fffb19ffe83c;
assign w_fix[98]='h000097ffe582fffa4b00071dfff580;
assign w_fix[99]='hfffc4a0006de0009f1fff4bf00189a;
assign w_fix[100]='hffffdd000a01000852fffbc60010e5;
assign w_fix[101]='hfffe12fff6ac000dc900012bfffc9d;
assign w_fix[102]='h00000d000f2a0005bb00050f001543;
assign w_fix[103]='hfff408fff6aa000818001f10ffe8f9;
assign w_fix[104]='hffff15ffff87000248fffe36000eea;
assign w_fix[105]='h00017b00141c0019930008c30019f0;
assign w_fix[106]='h00077a0010a70000ba000b40fffabf;
assign w_fix[107]='hffffa3000719fff40bfff422fffb6c;
assign w_fix[108]='hfff56c000a02000112000530fff20c;
assign w_fix[109]='h000107000fea00087c00099d0014e1;
assign w_fix[110]='h000a47fff33500053effd082000e36;
assign w_fix[111]='hfff7eb0007f6000cad00081ffffb30;
assign w_fix[112]='h00104c00014dfffaa5ffe9aa003f1d;
assign w_fix[113]='h00050e00076d000a27ffe70f0023bf;
assign w_fix[114]='hffff4effec0efff951ffdbb5fffc02;
assign w_fix[115]='h0002edfff6a0ffdeaafff953ffdfc7;
assign w_fix[116]='h00006100135600072d0009ca000f76;
assign w_fix[117]='hfff3abffff71fffbd900164bfff2e9;
assign w_fix[118]='h0001e2000892000c46ffeb6c00273e;
assign w_fix[119]='h000086fffc4d00003dfffe4e000510;
assign w_fix[120]='h0011c7ffeab2ffd4cf001d3effffdc;
assign w_fix[121]='hfffc2f001cb3fff7e9ffe8b0001094;
assign w_fix[122]='hfff68efffffeffeec40002affff93e;
assign w_fix[123]='h0002ab0008adffc600001545fff60e;
assign w_fix[124]='h0000c400054cffe91d0001e10012eb;
assign w_fix[125]='hfffce3000883ffc7c9ffe7740006e3;
assign w_fix[126]='h00036c000bc6ffc4f80006b8fffabc;
assign w_fix[127]='h00014700064900328d00088ffffb16;
assign w_fix[128]='h000730ffff57fffcb7ffef43000912;
assign w_fix[129]='hfff76ffff91800169f000574fff75b;
assign w_fix[130]='hfffeb7fffddaffff66fffcf10003c5;
assign w_fix[131]='h00023800050cffcf40000d58fff7f7;
assign w_fix[132]='hfffd64fffca5fff0cbffffa6000165;
assign w_fix[133]='hfff3c40013a6004b94fffb910004e6;
assign w_fix[134]='hfffeda000031fffb27fff819fffd38;
assign w_fix[135]='h0007f500038a00412f000ce90003eb;
assign w_fix[136]='h000986001c54000c910019f2fff2e4;
assign w_fix[137]='hfffadf0004d8ffe6bdffe8fd00035f;
assign w_fix[138]='h000034fffd5b004644fffe6bfff82f;
assign w_fix[139]='hffffeefff98100078bfffc8a0011cd;
assign w_fix[140]='h0006d0fff6c5ffbe40fffc8cfffadd;
assign w_fix[141]='hfff77a000622fff95100007afff7a3;
assign w_fix[142]='h000d1c000212ffe33000043c00017d;
assign w_fix[143]='hfffc09fff5e7ffdc3bfff4ba0001f7;
assign w_fix[144]='hffff260003b1fffe320001a0fff928;
assign w_fix[145]='hfffe73ffe9ebfffa72000d81ffe89e;
assign w_fix[146]='h00032dfffe34fffe4d000dc00007ad;
assign w_fix[147]='hfffd7cffff38004799fffb2b000a05;
assign w_fix[148]='h0000a7fffcaffff743fffa1c000326;
assign w_fix[149]='h0000c80001070005bb0004d2fffccb;
assign w_fix[150]='hfffc750002a2000a31fff6ccfffb28;
assign w_fix[151]='h0000ca00088a000309000e5ffff337;
assign w_fix[152]='hfffe7b0008d2fffb18000208fff878;
assign w_fix[153]='hffff3e000b1fffe9cdfffc97000a95;
assign w_fix[154]='h00003b000268000eb4fffcd3ffe9da;
assign w_fix[155]='hffff08000439ffe7b1000053000906;
assign w_fix[156]='hfffaa4000362ffe9720011defffd78;
assign w_fix[157]='h0000fd0002f2ffff16fffd100005a9;
assign w_fix[158]='hffffee00017affdce50000c7000258;
assign w_fix[159]='h000139fffd99000b11000218fff46b;
assign w_fix[160]='h000043fffdb60005ceffff5ffff5fa;
assign w_fix[161]='hffff110008d5fff380fffe28fffa8e;
assign w_fix[162]='h00013b0000e300070b00068bffed4c;
assign w_fix[163]='h0006da00099d000f18fff3b4000e5d;
assign w_fix[164]='hffffab0000bdfffdf2000337000376;
assign w_fix[165]='h0003080006e4001f23fffdb0fffb6b;
assign w_fix[166]='h0001fc001cc0000811000150fff8c9;
assign w_fix[167]='hfffd6e00044600032600049b000789;
assign w_fix[168]='h0001290005d9000961fffb78fffb15;
assign w_fix[169]='hffff5efffc760016d30000c4fffea8;
assign w_fix[170]='h0000b7fffd80001875fffa4fffec28;
assign w_fix[171]='hffff04000ddf0013aafff957ffea06;
assign w_fix[172]='hfff95c000ba0fff418000e2ffffa16;
assign w_fix[173]='h000013fff48a0001a2000f08ffedd3;
assign w_fix[174]='hfffe430007c0ffe383fff870ffffa9;
assign w_fix[175]='hffff0ffff407fff994fff65d00107d;
assign w_fix[176]='h0000a90001d7000da30003b5000173;
assign w_fix[177]='h0001c0ffff42fffcd0fff586000541;
assign w_fix[178]='h000096fffcc10002e5000a3efff347;
assign w_fix[179]='h00002c0000a2fff93200023b000a11;

endmodule