module createAandB_sigmoid #(
parameter aDW = 18,
parameter bDW = 18,
parameter numOfDots = 391, //�����зֵ�ĸ������������Ҷ˵�
parameter MW = 9
)(
input wire en,
input wire rst_n,
input wire [MW : 0] i,
output reg [(aDW - 1) : 0] a,
output reg [(bDW - 1) : 0] b
);

wire EN;

wire [(aDW - 1) : 0] aList [(numOfDots - 1) : 0];
wire [(bDW - 1) : 0] bList [(numOfDots - 1) : 0];

// assign aList[0] = 16'h0000; 
// assign aList[1] = 16'h0023; 
// assign aList[2] = 16'h008a; 
// assign aList[3] = 16'h0119; 
// assign aList[4] = 16'h01cb; 
// assign aList[5] = 16'h02e6; 
// assign aList[6] = 16'h041a; 
// assign aList[7] = 16'h052c; 
// assign aList[8] = 16'h067b; 
// assign aList[9] = 16'h0813; 
// assign aList[10] = 16'h09fb; 
// assign aList[11] = 16'h0c37; 
// assign aList[12] = 16'h0ec5; 
// assign aList[13] = 16'h119a; 
// assign aList[14] = 16'h149f; 
// assign aList[15] = 16'h17ad; 
// assign aList[16] = 16'h1a90; 
// assign aList[17] = 16'h1d0a; 
// assign aList[18] = 16'h1edd; 
// assign aList[19] = 16'h1fd6; 
// assign aList[20] = 16'h1fd6; 
// assign aList[21] = 16'h1edd; 
// assign aList[22] = 16'h1d0a; 
// assign aList[23] = 16'h1a90; 
// assign aList[24] = 16'h17ad; 
// assign aList[25] = 16'h149f; 
// assign aList[26] = 16'h119a; 
// assign aList[27] = 16'h0ec5; 
// assign aList[28] = 16'h0c37; 
// assign aList[29] = 16'h09fb; 
// assign aList[30] = 16'h0813; 
// assign aList[31] = 16'h067b; 
// assign aList[32] = 16'h052c; 
// assign aList[33] = 16'h041a; 
// assign aList[34] = 16'h02e6; 
// assign aList[35] = 16'h01cb; 
// assign aList[36] = 16'h0119; 
// assign aList[37] = 16'h008a; 
// assign aList[38] = 16'h0023; 

// assign bList[0] = 16'h0000;
// assign bList[1] = 16'h0123;
// assign bList[2] = 16'h038f;
// assign bList[3] = 16'h065a;
// assign bList[4] = 16'h0978;
// assign bList[5] = 16'h0de6;
// assign bList[6] = 16'h121d;
// assign bList[7] = 16'h1595;
// assign bList[8] = 16'h1984;
// assign bList[9] = 16'h1de6;
// assign bList[10] =16'h22a9;
// assign bList[11] = 16'h27af;
// assign bList[12] = 16'h2ccb;
// assign bList[13] = 16'h31c1;
// assign bList[14] = 16'h3648;
// assign bList[15] = 16'h3a1a;
// assign bList[16] = 16'h3cfd;
// assign bList[17] = 16'h3ed8;
// assign bList[18] = 16'h3fc2;
// assign bList[19] = 16'h4000;
// assign bList[20] = 16'h4000;
// assign bList[21] = 16'h403e;
// assign bList[22] = 16'h4128;
// assign bList[23] = 16'h4303;
// assign bList[24] = 16'h45e6;
// assign bList[25] = 16'h49b8;
// assign bList[26] = 16'h4e3f;
// assign bList[27] = 16'h5335;
// assign bList[28] = 16'h5851;
// assign bList[29] = 16'h5d57;
// assign bList[30] = 16'h621a;
// assign bList[31] = 16'h667c;
// assign bList[32] = 16'h6a6b;
// assign bList[33] = 16'h6de3;
// assign bList[34] = 16'h721a;
// assign bList[35] = 16'h7688;
// assign bList[36] = 16'h79a6;
// assign bList[37] = 16'h7c71;
// assign bList[38] = 16'h7edd;

assign aList[0] = 18'h00000; 
assign aList[1] = 18'h00032; 
assign aList[2] = 18'h00040; 
assign aList[3] = 18'h00052; 
assign aList[4] = 18'h0006a; 
assign aList[5] = 18'h00088; 
assign aList[6] = 18'h000a3; 
assign aList[7] = 18'h000b9; 
assign aList[8] = 18'h000d1; 
assign aList[9] = 18'h000ed; 
assign aList[10] = 18'h0010c; 
assign aList[11] = 18'h00130; 
assign aList[12] = 18'h00158; 
assign aList[13] = 18'h00186; 
assign aList[14] = 18'h001b9; 
assign aList[15] = 18'h001f4; 
assign aList[16] = 18'h00236; 
assign aList[17] = 18'h00280; 
assign aList[18] = 18'h002be; 
assign aList[19] = 18'h002eb; 
assign aList[20] = 18'h0031a; 
assign aList[21] = 18'h0034d; 
assign aList[22] = 18'h00383; 
assign aList[23] = 18'h003bc; 
assign aList[24] = 18'h003f9; 
assign aList[25] = 18'h00439; 
assign aList[26] = 18'h0047e; 
assign aList[27] = 18'h004c6; 
assign aList[28] = 18'h00514; 
assign aList[29] = 18'h00566; 
assign aList[30] = 18'h005bd; 
assign aList[31] = 18'h00619; 
assign aList[32] = 18'h0067b; 
assign aList[33] = 18'h006e3; 
assign aList[34] = 18'h00752; 
assign aList[35] = 18'h007c7; 
assign aList[36] = 18'h00843; 
assign aList[37] = 18'h008c7; 
assign aList[38] = 18'h00952; 
assign aList[39] = 18'h009e6; 
assign aList[40] = 18'h00a83; 
assign aList[41] = 18'h00afe; 
assign aList[42] = 18'h00b53; 
assign aList[43] = 18'h00bab; 
assign aList[44] = 18'h00c05; 
assign aList[45] = 18'h00c62; 
assign aList[46] = 18'h00cc1; 
assign aList[47] = 18'h00d24; 
assign aList[48] = 18'h00d88; 
assign aList[49] = 18'h00df0; 
assign aList[50] = 18'h00e5b; 
assign aList[51] = 18'h00ec9; 
assign aList[52] = 18'h00f3a; 
assign aList[53] = 18'h00fad; 
assign aList[54] = 18'h01025; 
assign aList[55] = 18'h0109f; 
assign aList[56] = 18'h0111d; 
assign aList[57] = 18'h0119e; 
assign aList[58] = 18'h01222; 
assign aList[59] = 18'h012ab; 
assign aList[60] = 18'h01336; 
assign aList[61] = 18'h013c6; 
assign aList[62] = 18'h01459; 
assign aList[63] = 18'h014f1; 
assign aList[64] = 18'h0158c; 
assign aList[65] = 18'h0162b; 
assign aList[66] = 18'h016ce; 
assign aList[67] = 18'h01776; 
assign aList[68] = 18'h01822; 
assign aList[69] = 18'h018d2; 
assign aList[70] = 18'h01986; 
assign aList[71] = 18'h01a3f; 
assign aList[72] = 18'h01afd; 
assign aList[73] = 18'h01bbf; 
assign aList[74] = 18'h01c85; 
assign aList[75] = 18'h01d51; 
assign aList[76] = 18'h01e21; 
assign aList[77] = 18'h01ef7; 
assign aList[78] = 18'h01fd1; 
assign aList[79] = 18'h020b0; 
assign aList[80] = 18'h02194; 
assign aList[81] = 18'h0227d; 
assign aList[82] = 18'h0236c; 
assign aList[83] = 18'h0245f; 
assign aList[84] = 18'h02558; 
assign aList[85] = 18'h02656; 
assign aList[86] = 18'h02759; 
assign aList[87] = 18'h02862; 
assign aList[88] = 18'h02970; 
assign aList[89] = 18'h02a83; 
assign aList[90] = 18'h02b9c; 
assign aList[91] = 18'h02cba; 
assign aList[92] = 18'h02ddd; 
assign aList[93] = 18'h02f06; 
assign aList[94] = 18'h03034; 
assign aList[95] = 18'h03167; 
assign aList[96] = 18'h0329f; 
assign aList[97] = 18'h033dc; 
assign aList[98] = 18'h0351f; 
assign aList[99] = 18'h03666; 
assign aList[100] = 18'h037b3; 
assign aList[101] = 18'h038af; 
assign aList[102] = 18'h03959; 
assign aList[103] = 18'h03a04; 
assign aList[104] = 18'h03ab0; 
assign aList[105] = 18'h03b5d; 
assign aList[106] = 18'h03c0c; 
assign aList[107] = 18'h03cbb; 
assign aList[108] = 18'h03d6c; 
assign aList[109] = 18'h03e1e; 
assign aList[110] = 18'h03ed1; 
assign aList[111] = 18'h03f84; 
assign aList[112] = 18'h04039; 
assign aList[113] = 18'h040ef; 
assign aList[114] = 18'h041a6; 
assign aList[115] = 18'h0425e; 
assign aList[116] = 18'h04316; 
assign aList[117] = 18'h043d0; 
assign aList[118] = 18'h0448a; 
assign aList[119] = 18'h04546; 
assign aList[120] = 18'h04602; 
assign aList[121] = 18'h046bf; 
assign aList[122] = 18'h0477c; 
assign aList[123] = 18'h0483b; 
assign aList[124] = 18'h048fa; 
assign aList[125] = 18'h049b9; 
assign aList[126] = 18'h04a7a; 
assign aList[127] = 18'h04b3b; 
assign aList[128] = 18'h04bfc; 
assign aList[129] = 18'h04cbe; 
assign aList[130] = 18'h04d80; 
assign aList[131] = 18'h04e43; 
assign aList[132] = 18'h04f07; 
assign aList[133] = 18'h04fca; 
assign aList[134] = 18'h0508e; 
assign aList[135] = 18'h05153; 
assign aList[136] = 18'h05217; 
assign aList[137] = 18'h052dc; 
assign aList[138] = 18'h053a1; 
assign aList[139] = 18'h05466; 
assign aList[140] = 18'h0552b; 
assign aList[141] = 18'h055f0; 
assign aList[142] = 18'h056b5; 
assign aList[143] = 18'h0577a; 
assign aList[144] = 18'h0583f; 
assign aList[145] = 18'h05903; 
assign aList[146] = 18'h059c8; 
assign aList[147] = 18'h05a8c; 
assign aList[148] = 18'h05b50; 
assign aList[149] = 18'h05c13; 
assign aList[150] = 18'h05cd6; 
assign aList[151] = 18'h05d98; 
assign aList[152] = 18'h05e5a; 
assign aList[153] = 18'h05f1b; 
assign aList[154] = 18'h05fdc; 
assign aList[155] = 18'h0609b; 
assign aList[156] = 18'h0615a; 
assign aList[157] = 18'h06219; 
assign aList[158] = 18'h062d6; 
assign aList[159] = 18'h06392; 
assign aList[160] = 18'h0644d; 
assign aList[161] = 18'h06507; 
assign aList[162] = 18'h065c0; 
assign aList[163] = 18'h06678; 
assign aList[164] = 18'h0672e; 
assign aList[165] = 18'h067e3; 
assign aList[166] = 18'h06897; 
assign aList[167] = 18'h06949; 
assign aList[168] = 18'h069fa; 
assign aList[169] = 18'h06aa9; 
assign aList[170] = 18'h06b56; 
assign aList[171] = 18'h06c02; 
assign aList[172] = 18'h06cab; 
assign aList[173] = 18'h06da6; 
assign aList[174] = 18'h06eef; 
assign aList[175] = 18'h0702e; 
assign aList[176] = 18'h07165; 
assign aList[177] = 18'h07293; 
assign aList[178] = 18'h073b7; 
assign aList[179] = 18'h074d0; 
assign aList[180] = 18'h075df; 
assign aList[181] = 18'h076e3; 
assign aList[182] = 18'h077da; 
assign aList[183] = 18'h078c6; 
assign aList[184] = 18'h079a5; 
assign aList[185] = 18'h07a78; 
assign aList[186] = 18'h07b3d; 
assign aList[187] = 18'h07bf4; 
assign aList[188] = 18'h07c9d; 
assign aList[189] = 18'h07d38; 
assign aList[190] = 18'h07dc4; 
assign aList[191] = 18'h07e41; 
assign aList[192] = 18'h07eb0; 
assign aList[193] = 18'h07f36; 
assign aList[194] = 18'h07fb5; 
assign aList[195] = 18'h07ff5; 
assign aList[196] = 18'h07ff5; 
assign aList[197] = 18'h07fb5; 
assign aList[198] = 18'h07f36; 
assign aList[199] = 18'h07eb0; 
assign aList[200] = 18'h07e41; 
assign aList[201] = 18'h07dc4; 
assign aList[202] = 18'h07d38; 
assign aList[203] = 18'h07c9d; 
assign aList[204] = 18'h07bf4; 
assign aList[205] = 18'h07b3d; 
assign aList[206] = 18'h07a78; 
assign aList[207] = 18'h079a5; 
assign aList[208] = 18'h078c6; 
assign aList[209] = 18'h077da; 
assign aList[210] = 18'h076e3; 
assign aList[211] = 18'h075df; 
assign aList[212] = 18'h074d0; 
assign aList[213] = 18'h073b7; 
assign aList[214] = 18'h07293; 
assign aList[215] = 18'h07165; 
assign aList[216] = 18'h0702e; 
assign aList[217] = 18'h06eef; 
assign aList[218] = 18'h06da6; 
assign aList[219] = 18'h06cab; 
assign aList[220] = 18'h06c02; 
assign aList[221] = 18'h06b56; 
assign aList[222] = 18'h06aa9; 
assign aList[223] = 18'h069fa; 
assign aList[224] = 18'h06949; 
assign aList[225] = 18'h06897; 
assign aList[226] = 18'h067e3; 
assign aList[227] = 18'h0672e; 
assign aList[228] = 18'h06678; 
assign aList[229] = 18'h065c0; 
assign aList[230] = 18'h06507; 
assign aList[231] = 18'h0644d; 
assign aList[232] = 18'h06392; 
assign aList[233] = 18'h062d6; 
assign aList[234] = 18'h06219; 
assign aList[235] = 18'h0615a; 
assign aList[236] = 18'h0609b; 
assign aList[237] = 18'h05fdc; 
assign aList[238] = 18'h05f1b; 
assign aList[239] = 18'h05e5a; 
assign aList[240] = 18'h05d98; 
assign aList[241] = 18'h05cd6; 
assign aList[242] = 18'h05c13; 
assign aList[243] = 18'h05b50; 
assign aList[244] = 18'h05a8c; 
assign aList[245] = 18'h059c8; 
assign aList[246] = 18'h05903; 
assign aList[247] = 18'h0583f; 
assign aList[248] = 18'h0577a; 
assign aList[249] = 18'h056b5; 
assign aList[250] = 18'h055f0; 
assign aList[251] = 18'h0552b; 
assign aList[252] = 18'h05466; 
assign aList[253] = 18'h053a1; 
assign aList[254] = 18'h052dc; 
assign aList[255] = 18'h05217; 
assign aList[256] = 18'h05153; 
assign aList[257] = 18'h0508e; 
assign aList[258] = 18'h04fca; 
assign aList[259] = 18'h04f07; 
assign aList[260] = 18'h04e43; 
assign aList[261] = 18'h04d80; 
assign aList[262] = 18'h04cbe; 
assign aList[263] = 18'h04bfc; 
assign aList[264] = 18'h04b3b; 
assign aList[265] = 18'h04a7a; 
assign aList[266] = 18'h049b9; 
assign aList[267] = 18'h048fa; 
assign aList[268] = 18'h0483b; 
assign aList[269] = 18'h0477c; 
assign aList[270] = 18'h046bf; 
assign aList[271] = 18'h04602; 
assign aList[272] = 18'h04546; 
assign aList[273] = 18'h0448a; 
assign aList[274] = 18'h043d0; 
assign aList[275] = 18'h04316; 
assign aList[276] = 18'h0425e; 
assign aList[277] = 18'h041a6; 
assign aList[278] = 18'h040ef; 
assign aList[279] = 18'h04039; 
assign aList[280] = 18'h03f84; 
assign aList[281] = 18'h03ed1; 
assign aList[282] = 18'h03e1e; 
assign aList[283] = 18'h03d6c; 
assign aList[284] = 18'h03cbb; 
assign aList[285] = 18'h03c0c; 
assign aList[286] = 18'h03b5d; 
assign aList[287] = 18'h03ab0; 
assign aList[288] = 18'h03a04; 
assign aList[289] = 18'h03959; 
assign aList[290] = 18'h038af; 
assign aList[291] = 18'h037b3; 
assign aList[292] = 18'h03666; 
assign aList[293] = 18'h0351f; 
assign aList[294] = 18'h033dc; 
assign aList[295] = 18'h0329f; 
assign aList[296] = 18'h03167; 
assign aList[297] = 18'h03034; 
assign aList[298] = 18'h02f06; 
assign aList[299] = 18'h02ddd; 
assign aList[300] = 18'h02cba; 
assign aList[301] = 18'h02b9c; 
assign aList[302] = 18'h02a83; 
assign aList[303] = 18'h02970; 
assign aList[304] = 18'h02862; 
assign aList[305] = 18'h02759; 
assign aList[306] = 18'h02656; 
assign aList[307] = 18'h02558; 
assign aList[308] = 18'h0245f; 
assign aList[309] = 18'h0236c; 
assign aList[310] = 18'h0227d; 
assign aList[311] = 18'h02194; 
assign aList[312] = 18'h020b0; 
assign aList[313] = 18'h01fd1; 
assign aList[314] = 18'h01ef7; 
assign aList[315] = 18'h01e21; 
assign aList[316] = 18'h01d51; 
assign aList[317] = 18'h01c85; 
assign aList[318] = 18'h01bbf; 
assign aList[319] = 18'h01afd; 
assign aList[320] = 18'h01a3f; 
assign aList[321] = 18'h01986; 
assign aList[322] = 18'h018d2; 
assign aList[323] = 18'h01822; 
assign aList[324] = 18'h01776; 
assign aList[325] = 18'h016ce; 
assign aList[326] = 18'h0162b; 
assign aList[327] = 18'h0158c; 
assign aList[328] = 18'h014f1; 
assign aList[329] = 18'h01459; 
assign aList[330] = 18'h013c6; 
assign aList[331] = 18'h01336; 
assign aList[332] = 18'h012ab; 
assign aList[333] = 18'h01222; 
assign aList[334] = 18'h0119e; 
assign aList[335] = 18'h0111d; 
assign aList[336] = 18'h0109f; 
assign aList[337] = 18'h01025; 
assign aList[338] = 18'h00fad; 
assign aList[339] = 18'h00f3a; 
assign aList[340] = 18'h00ec9; 
assign aList[341] = 18'h00e5b; 
assign aList[342] = 18'h00df0; 
assign aList[343] = 18'h00d88; 
assign aList[344] = 18'h00d24; 
assign aList[345] = 18'h00cc1; 
assign aList[346] = 18'h00c62; 
assign aList[347] = 18'h00c05; 
assign aList[348] = 18'h00bab; 
assign aList[349] = 18'h00b53; 
assign aList[350] = 18'h00afe; 
assign aList[351] = 18'h00a83; 
assign aList[352] = 18'h009e6; 
assign aList[353] = 18'h00952; 
assign aList[354] = 18'h008c7; 
assign aList[355] = 18'h00843; 
assign aList[356] = 18'h007c7; 
assign aList[357] = 18'h00752; 
assign aList[358] = 18'h006e3; 
assign aList[359] = 18'h0067b; 
assign aList[360] = 18'h00619; 
assign aList[361] = 18'h005bd; 
assign aList[362] = 18'h00566; 
assign aList[363] = 18'h00514; 
assign aList[364] = 18'h004c6; 
assign aList[365] = 18'h0047e; 
assign aList[366] = 18'h00439; 
assign aList[367] = 18'h003f9; 
assign aList[368] = 18'h003bc; 
assign aList[369] = 18'h00383; 
assign aList[370] = 18'h0034d; 
assign aList[371] = 18'h0031a; 
assign aList[372] = 18'h002eb; 
assign aList[373] = 18'h002be; 
assign aList[374] = 18'h00280; 
assign aList[375] = 18'h00236; 
assign aList[376] = 18'h001f4; 
assign aList[377] = 18'h001b9; 
assign aList[378] = 18'h00186; 
assign aList[379] = 18'h00158; 
assign aList[380] = 18'h00130; 
assign aList[381] = 18'h0010c; 
assign aList[382] = 18'h000ed; 
assign aList[383] = 18'h000d1; 
assign aList[384] = 18'h000b9; 
assign aList[385] = 18'h000a3; 
assign aList[386] = 18'h00088; 
assign aList[387] = 18'h0006a; 
assign aList[388] = 18'h00052; 
assign aList[389] = 18'h00040; 
assign aList[390] = 18'h00032; 

assign bList[0] = 18'h00000; 
assign bList[1] = 18'h001bb; 
assign bList[2] = 18'h00229; 
assign bList[3] = 18'h002b1; 
assign bList[4] = 18'h0035a; 
assign bList[5] = 18'h0042c; 
assign bList[6] = 18'h004e6; 
assign bList[7] = 18'h00575; 
assign bList[8] = 18'h00615; 
assign bList[9] = 18'h006c6; 
assign bList[10] = 18'h0078a; 
assign bList[11] = 18'h00864; 
assign bList[12] = 18'h00956; 
assign bList[13] = 18'h00a61; 
assign bList[14] = 18'h00b8a; 
assign bList[15] = 18'h00cd2; 
assign bList[16] = 18'h00e3c; 
assign bList[17] = 18'h00fcd; 
assign bList[18] = 18'h01112; 
assign bList[19] = 18'h011fb; 
assign bList[20] = 18'h012ee; 
assign bList[21] = 18'h013ee; 
assign bList[22] = 18'h014fb; 
assign bList[23] = 18'h01615; 
assign bList[24] = 18'h0173d; 
assign bList[25] = 18'h01873; 
assign bList[26] = 18'h019b9; 
assign bList[27] = 18'h01b0e; 
assign bList[28] = 18'h01c73; 
assign bList[29] = 18'h01de9; 
assign bList[30] = 18'h01f71; 
assign bList[31] = 18'h0210b; 
assign bList[32] = 18'h022b8; 
assign bList[33] = 18'h02479; 
assign bList[34] = 18'h0264f; 
assign bList[35] = 18'h02839; 
assign bList[36] = 18'h02a39; 
assign bList[37] = 18'h02c50; 
assign bList[38] = 18'h02e7e; 
assign bList[39] = 18'h030c4; 
assign bList[40] = 18'h03323; 
assign bList[41] = 18'h034f9; 
assign bList[42] = 18'h0363b; 
assign bList[43] = 18'h03784; 
assign bList[44] = 18'h038d4; 
assign bList[45] = 18'h03a2a; 
assign bList[46] = 18'h03b87; 
assign bList[47] = 18'h03ceb; 
assign bList[48] = 18'h03e56; 
assign bList[49] = 18'h03fc8; 
assign bList[50] = 18'h04141; 
assign bList[51] = 18'h042c1; 
assign bList[52] = 18'h04448; 
assign bList[53] = 18'h045d6; 
assign bList[54] = 18'h0476c; 
assign bList[55] = 18'h04909; 
assign bList[56] = 18'h04aad; 
assign bList[57] = 18'h04c59; 
assign bList[58] = 18'h04e0c; 
assign bList[59] = 18'h04fc7; 
assign bList[60] = 18'h05189; 
assign bList[61] = 18'h05353; 
assign bList[62] = 18'h05524; 
assign bList[63] = 18'h056fc; 
assign bList[64] = 18'h058dd; 
assign bList[65] = 18'h05ac4; 
assign bList[66] = 18'h05cb3; 
assign bList[67] = 18'h05eaa; 
assign bList[68] = 18'h060a8; 
assign bList[69] = 18'h062ad; 
assign bList[70] = 18'h064b9; 
assign bList[71] = 18'h066cd; 
assign bList[72] = 18'h068e8; 
assign bList[73] = 18'h06b0a; 
assign bList[74] = 18'h06d33; 
assign bList[75] = 18'h06f62; 
assign bList[76] = 18'h07199; 
assign bList[77] = 18'h073d6; 
assign bList[78] = 18'h07619; 
assign bList[79] = 18'h07863; 
assign bList[80] = 18'h07ab3; 
assign bList[81] = 18'h07d09; 
assign bList[82] = 18'h07f64; 
assign bList[83] = 18'h081c5; 
assign bList[84] = 18'h0842b; 
assign bList[85] = 18'h08697; 
assign bList[86] = 18'h08907; 
assign bList[87] = 18'h08b7b; 
assign bList[88] = 18'h08df4; 
assign bList[89] = 18'h09070; 
assign bList[90] = 18'h092f0; 
assign bList[91] = 18'h09574; 
assign bList[92] = 18'h097fa; 
assign bList[93] = 18'h09a83; 
assign bList[94] = 18'h09d0e; 
assign bList[95] = 18'h09f9a; 
assign bList[96] = 18'h0a228; 
assign bList[97] = 18'h0a4b7; 
assign bList[98] = 18'h0a746; 
assign bList[99] = 18'h0a9d5; 
assign bList[100] = 18'h0ac63; 
assign bList[101] = 18'h0ae4c; 
assign bList[102] = 18'h0af93; 
assign bList[103] = 18'h0b0d9; 
assign bList[104] = 18'h0b21e; 
assign bList[105] = 18'h0b363; 
assign bList[106] = 18'h0b4a7; 
assign bList[107] = 18'h0b5eb; 
assign bList[108] = 18'h0b72e; 
assign bList[109] = 18'h0b870; 
assign bList[110] = 18'h0b9b1; 
assign bList[111] = 18'h0baf2; 
assign bList[112] = 18'h0bc31; 
assign bList[113] = 18'h0bd6f; 
assign bList[114] = 18'h0beac; 
assign bList[115] = 18'h0bfe8; 
assign bList[116] = 18'h0c123; 
assign bList[117] = 18'h0c25c; 
assign bList[118] = 18'h0c393; 
assign bList[119] = 18'h0c4ca; 
assign bList[120] = 18'h0c5fe; 
assign bList[121] = 18'h0c731; 
assign bList[122] = 18'h0c862; 
assign bList[123] = 18'h0c992; 
assign bList[124] = 18'h0cabf; 
assign bList[125] = 18'h0cbeb; 
assign bList[126] = 18'h0cd14; 
assign bList[127] = 18'h0ce3c; 
assign bList[128] = 18'h0cf61; 
assign bList[129] = 18'h0d084; 
assign bList[130] = 18'h0d1a5; 
assign bList[131] = 18'h0d2c3; 
assign bList[132] = 18'h0d3df; 
assign bList[133] = 18'h0d4f8; 
assign bList[134] = 18'h0d60f; 
assign bList[135] = 18'h0d723; 
assign bList[136] = 18'h0d834; 
assign bList[137] = 18'h0d943; 
assign bList[138] = 18'h0da4e; 
assign bList[139] = 18'h0db57; 
assign bList[140] = 18'h0dc5d; 
assign bList[141] = 18'h0dd5f; 
assign bList[142] = 18'h0de5f; 
assign bList[143] = 18'h0df5b; 
assign bList[144] = 18'h0e054; 
assign bList[145] = 18'h0e14a; 
assign bList[146] = 18'h0e23c; 
assign bList[147] = 18'h0e32b; 
assign bList[148] = 18'h0e417; 
assign bList[149] = 18'h0e4ff; 
assign bList[150] = 18'h0e5e3; 
assign bList[151] = 18'h0e6c4; 
assign bList[152] = 18'h0e7a1; 
assign bList[153] = 18'h0e87a; 
assign bList[154] = 18'h0e950; 
assign bList[155] = 18'h0ea22; 
assign bList[156] = 18'h0eaf0; 
assign bList[157] = 18'h0ebba; 
assign bList[158] = 18'h0ec80; 
assign bList[159] = 18'h0ed42; 
assign bList[160] = 18'h0ee00; 
assign bList[161] = 18'h0eeba; 
assign bList[162] = 18'h0ef70; 
assign bList[163] = 18'h0f022; 
assign bList[164] = 18'h0f0d0; 
assign bList[165] = 18'h0f179; 
assign bList[166] = 18'h0f21f; 
assign bList[167] = 18'h0f2c0; 
assign bList[168] = 18'h0f35e; 
assign bList[169] = 18'h0f3f7; 
assign bList[170] = 18'h0f48c; 
assign bList[171] = 18'h0f51d; 
assign bList[172] = 18'h0f5a9; 
assign bList[173] = 18'h0f675; 
assign bList[174] = 18'h0f776; 
assign bList[175] = 18'h0f865; 
assign bList[176] = 18'h0f945; 
assign bList[177] = 18'h0fa14; 
assign bList[178] = 18'h0fad4; 
assign bList[179] = 18'h0fb84; 
assign bList[180] = 18'h0fc25; 
assign bList[181] = 18'h0fcb7; 
assign bList[182] = 18'h0fd3a; 
assign bList[183] = 18'h0fdb0; 
assign bList[184] = 18'h0fe19; 
assign bList[185] = 18'h0fe75; 
assign bList[186] = 18'h0fec5; 
assign bList[187] = 18'h0ff09; 
assign bList[188] = 18'h0ff44; 
assign bList[189] = 18'h0ff74; 
assign bList[190] = 18'h0ff9b; 
assign bList[191] = 18'h0ffbb; 
assign bList[192] = 18'h0ffd3; 
assign bList[193] = 18'h0ffec; 
assign bList[194] = 18'h0fffc; 
assign bList[195] = 18'h10000; 
assign bList[196] = 18'h10000; 
assign bList[197] = 18'h10004; 
assign bList[198] = 18'h10014; 
assign bList[199] = 18'h1002d; 
assign bList[200] = 18'h10045; 
assign bList[201] = 18'h10065; 
assign bList[202] = 18'h1008c; 
assign bList[203] = 18'h100bc; 
assign bList[204] = 18'h100f7; 
assign bList[205] = 18'h1013b; 
assign bList[206] = 18'h1018b; 
assign bList[207] = 18'h101e7; 
assign bList[208] = 18'h10250; 
assign bList[209] = 18'h102c6; 
assign bList[210] = 18'h10349; 
assign bList[211] = 18'h103db; 
assign bList[212] = 18'h1047c; 
assign bList[213] = 18'h1052c; 
assign bList[214] = 18'h105ec; 
assign bList[215] = 18'h106bb; 
assign bList[216] = 18'h1079b; 
assign bList[217] = 18'h1088a; 
assign bList[218] = 18'h1098b; 
assign bList[219] = 18'h10a57; 
assign bList[220] = 18'h10ae3; 
assign bList[221] = 18'h10b74; 
assign bList[222] = 18'h10c09; 
assign bList[223] = 18'h10ca2; 
assign bList[224] = 18'h10d40; 
assign bList[225] = 18'h10de1; 
assign bList[226] = 18'h10e87; 
assign bList[227] = 18'h10f30; 
assign bList[228] = 18'h10fde; 
assign bList[229] = 18'h11090; 
assign bList[230] = 18'h11146; 
assign bList[231] = 18'h11200; 
assign bList[232] = 18'h112be; 
assign bList[233] = 18'h11380; 
assign bList[234] = 18'h11446; 
assign bList[235] = 18'h11510; 
assign bList[236] = 18'h115de; 
assign bList[237] = 18'h116b0; 
assign bList[238] = 18'h11786; 
assign bList[239] = 18'h1185f; 
assign bList[240] = 18'h1193c; 
assign bList[241] = 18'h11a1d; 
assign bList[242] = 18'h11b01; 
assign bList[243] = 18'h11be9; 
assign bList[244] = 18'h11cd5; 
assign bList[245] = 18'h11dc4; 
assign bList[246] = 18'h11eb6; 
assign bList[247] = 18'h11fac; 
assign bList[248] = 18'h120a5; 
assign bList[249] = 18'h121a1; 
assign bList[250] = 18'h122a1; 
assign bList[251] = 18'h123a3; 
assign bList[252] = 18'h124a9; 
assign bList[253] = 18'h125b2; 
assign bList[254] = 18'h126bd; 
assign bList[255] = 18'h127cc; 
assign bList[256] = 18'h128dd; 
assign bList[257] = 18'h129f1; 
assign bList[258] = 18'h12b08; 
assign bList[259] = 18'h12c21; 
assign bList[260] = 18'h12d3d; 
assign bList[261] = 18'h12e5b; 
assign bList[262] = 18'h12f7c; 
assign bList[263] = 18'h1309f; 
assign bList[264] = 18'h131c4; 
assign bList[265] = 18'h132ec; 
assign bList[266] = 18'h13415; 
assign bList[267] = 18'h13541; 
assign bList[268] = 18'h1366e; 
assign bList[269] = 18'h1379e; 
assign bList[270] = 18'h138cf; 
assign bList[271] = 18'h13a02; 
assign bList[272] = 18'h13b36; 
assign bList[273] = 18'h13c6d; 
assign bList[274] = 18'h13da4; 
assign bList[275] = 18'h13edd; 
assign bList[276] = 18'h14018; 
assign bList[277] = 18'h14154; 
assign bList[278] = 18'h14291; 
assign bList[279] = 18'h143cf; 
assign bList[280] = 18'h1450e; 
assign bList[281] = 18'h1464f; 
assign bList[282] = 18'h14790; 
assign bList[283] = 18'h148d2; 
assign bList[284] = 18'h14a15; 
assign bList[285] = 18'h14b59; 
assign bList[286] = 18'h14c9d; 
assign bList[287] = 18'h14de2; 
assign bList[288] = 18'h14f27; 
assign bList[289] = 18'h1506d; 
assign bList[290] = 18'h151b4; 
assign bList[291] = 18'h1539d; 
assign bList[292] = 18'h1562b; 
assign bList[293] = 18'h158ba; 
assign bList[294] = 18'h15b49; 
assign bList[295] = 18'h15dd8; 
assign bList[296] = 18'h16066; 
assign bList[297] = 18'h162f2; 
assign bList[298] = 18'h1657d; 
assign bList[299] = 18'h16806; 
assign bList[300] = 18'h16a8c; 
assign bList[301] = 18'h16d10; 
assign bList[302] = 18'h16f90; 
assign bList[303] = 18'h1720c; 
assign bList[304] = 18'h17485; 
assign bList[305] = 18'h176f9; 
assign bList[306] = 18'h17969; 
assign bList[307] = 18'h17bd5; 
assign bList[308] = 18'h17e3b; 
assign bList[309] = 18'h1809c; 
assign bList[310] = 18'h182f7; 
assign bList[311] = 18'h1854d; 
assign bList[312] = 18'h1879d; 
assign bList[313] = 18'h189e7; 
assign bList[314] = 18'h18c2a; 
assign bList[315] = 18'h18e67; 
assign bList[316] = 18'h1909e; 
assign bList[317] = 18'h192cd; 
assign bList[318] = 18'h194f6; 
assign bList[319] = 18'h19718; 
assign bList[320] = 18'h19933; 
assign bList[321] = 18'h19b47; 
assign bList[322] = 18'h19d53; 
assign bList[323] = 18'h19f58; 
assign bList[324] = 18'h1a156; 
assign bList[325] = 18'h1a34d; 
assign bList[326] = 18'h1a53c; 
assign bList[327] = 18'h1a723; 
assign bList[328] = 18'h1a904; 
assign bList[329] = 18'h1aadc; 
assign bList[330] = 18'h1acad; 
assign bList[331] = 18'h1ae77; 
assign bList[332] = 18'h1b039; 
assign bList[333] = 18'h1b1f4; 
assign bList[334] = 18'h1b3a7; 
assign bList[335] = 18'h1b553; 
assign bList[336] = 18'h1b6f7; 
assign bList[337] = 18'h1b894; 
assign bList[338] = 18'h1ba2a; 
assign bList[339] = 18'h1bbb8; 
assign bList[340] = 18'h1bd3f; 
assign bList[341] = 18'h1bebf; 
assign bList[342] = 18'h1c038; 
assign bList[343] = 18'h1c1aa; 
assign bList[344] = 18'h1c315; 
assign bList[345] = 18'h1c479; 
assign bList[346] = 18'h1c5d6; 
assign bList[347] = 18'h1c72c; 
assign bList[348] = 18'h1c87c; 
assign bList[349] = 18'h1c9c5; 
assign bList[350] = 18'h1cb07; 
assign bList[351] = 18'h1ccdd; 
assign bList[352] = 18'h1cf3c; 
assign bList[353] = 18'h1d182; 
assign bList[354] = 18'h1d3b0; 
assign bList[355] = 18'h1d5c7; 
assign bList[356] = 18'h1d7c7; 
assign bList[357] = 18'h1d9b1; 
assign bList[358] = 18'h1db87; 
assign bList[359] = 18'h1dd48; 
assign bList[360] = 18'h1def5; 
assign bList[361] = 18'h1e08f; 
assign bList[362] = 18'h1e217; 
assign bList[363] = 18'h1e38d; 
assign bList[364] = 18'h1e4f2; 
assign bList[365] = 18'h1e647; 
assign bList[366] = 18'h1e78d; 
assign bList[367] = 18'h1e8c3; 
assign bList[368] = 18'h1e9eb; 
assign bList[369] = 18'h1eb05; 
assign bList[370] = 18'h1ec12; 
assign bList[371] = 18'h1ed12; 
assign bList[372] = 18'h1ee05; 
assign bList[373] = 18'h1eeee; 
assign bList[374] = 18'h1f033; 
assign bList[375] = 18'h1f1c4; 
assign bList[376] = 18'h1f32e; 
assign bList[377] = 18'h1f476; 
assign bList[378] = 18'h1f59f; 
assign bList[379] = 18'h1f6aa; 
assign bList[380] = 18'h1f79c; 
assign bList[381] = 18'h1f876; 
assign bList[382] = 18'h1f93a; 
assign bList[383] = 18'h1f9eb; 
assign bList[384] = 18'h1fa8b; 
assign bList[385] = 18'h1fb1a; 
assign bList[386] = 18'h1fbd4; 
assign bList[387] = 18'h1fca6; 
assign bList[388] = 18'h1fd4f; 
assign bList[389] = 18'h1fdd7; 
assign bList[390] = 18'h1fe45; 

AND_2_1 AND_2_1_inst(
.IN_1   (   en      ),
.IN_0   (   rst_n   ),
.OUT    (   EN      )
);

always @* begin
    if(EN == 1'b1) begin
        a = aList[i];
    end
    else begin
        a = 'd0;
    end
end

always @* begin
    if(EN == 1'b1) begin
        b = bList[i];
    end
    else begin
        b = 'd0;
    end
end

endmodule
