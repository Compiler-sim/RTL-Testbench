module rf_buffer #(
  parameter D_WL = 24,
  parameter UNITS_NUM = 5
)(
   input [7:0] addr,
   output [UNITS_NUM*D_WL-1:0] w_o
);

wire [D_WL*UNITS_NUM-1:0] w_fix [0:179];
assign w_o = w_fix[addr];
assign w_fix[0]='h000045002207000cefffe393000b71;
assign w_fix[1]='hfff3b4fff724001a97ffebdcffef54;
assign w_fix[2]='hfff937000944001aadfff19dfff187;
assign w_fix[3]='hfffad3000973001560000140ffe816;
assign w_fix[4]='hfff9cd000f1a001415fff006fff8f3;
assign w_fix[5]='h00032c000f25001d89000893001c8c;
assign w_fix[6]='hfff84c001ee400106a000dcb00319b;
assign w_fix[7]='h00021dfffddcffef7400053600114d;
assign w_fix[8]='h0008c1fff810000be6001561fff544;
assign w_fix[9]='hffff55000566000e4fffffbbffe80f;
assign w_fix[10]='hffff74fffb2c000ac9fff89cffe85d;
assign w_fix[11]='h0002b60009f0000b95ffe021000d9d;
assign w_fix[12]='hfffd9b000554000ce7fff868ffeb7f;
assign w_fix[13]='h0006e7ffe6f4fff376fffee0fffa8d;
assign w_fix[14]='h000031fff2010009a00001c2ffee1a;
assign w_fix[15]='h0000befff07efff3e0fff114ffe875;
assign w_fix[16]='hfffc16001c9d0007a1ffef0effd961;
assign w_fix[17]='h00027800144e00102900010a000807;
assign w_fix[18]='hfffea4ffecf3fffff9fffa67fff30b;
assign w_fix[19]='h0000eafff9eafff8aefff4f2fff999;
assign w_fix[20]='hffffeffffb030000fc0005f3000e3b;
assign w_fix[21]='hfff09f00038d0012a1fff16a0009de;
assign w_fix[22]='hfff9000020ff0009a3000df8001856;
assign w_fix[23]='hfffe830009580013360000cfffda60;
assign w_fix[24]='hfffc50ffff1cfff7bb0000b5fff897;
assign w_fix[25]='h000be5000826ffe575001725001572;
assign w_fix[26]='hffff10000948fff166fffb94000477;
assign w_fix[27]='hfffc7bffe591fffaa6000887fff704;
assign w_fix[28]='hffff0afffabb000c590000fcffcffd;
assign w_fix[29]='h000307fffab7fff402000a35fffd21;
assign w_fix[30]='h001477ffe11dfffc4b0042fe002e99;
assign w_fix[31]='hfff8e6ffeed5fffd2d000028000123;
assign w_fix[32]='h0013c30011eefffe32000377000aef;
assign w_fix[33]='hffff2a0006560009eefff826fffd16;
assign w_fix[34]='h0000e1fffb2afffeb4fff6fafffabe;
assign w_fix[35]='hfffeb1fff3e3fffcfc0012c80009fe;
assign w_fix[36]='hfffcc8000241fffe75000e6b000e96;
assign w_fix[37]='hfffd79fff1f1000274fffbfbfff631;
assign w_fix[38]='hfff59a001280000e0a000e91fff630;
assign w_fix[39]='h000ab0fffe6ffffcf30004290002c5;
assign w_fix[40]='h00047ffff989fffd87ffff06000265;
assign w_fix[41]='h0016fa0007d40005d0000a0d0005cd;
assign w_fix[42]='h000fe0fffe8f0000acfff83d00030c;
assign w_fix[43]='hfff5a8000c6000024bffe4bdfff0ef;
assign w_fix[44]='h000008fff9c30000050007dc0006eb;
assign w_fix[45]='h00049efffaf0000430ffeba0fff5b4;
assign w_fix[46]='h001711fff03bfffcbfffe622fffe95;
assign w_fix[47]='h0004f5fffd9afffec3001135000e19;
assign w_fix[48]='h0003ed00005efffe55fff2dbfffbb3;
assign w_fix[49]='hffff4b0014de000088fff020fff5df;
assign w_fix[50]='h000eb9000016fff508003e56001187;
assign w_fix[51]='h001358fffb2afff72a00138600177d;
assign w_fix[52]='hffe9d90014460000e80018610011e6;
assign w_fix[53]='h000ddcfffa2100003d0002b5000426;
assign w_fix[54]='hfffc53ffe9e4fffe85000f02000ac5;
assign w_fix[55]='h0004f5000e26fffda20004cf00060e;
assign w_fix[56]='h00084dfff647fffe52fff752fffd9c;
assign w_fix[57]='hffecf10015a00000adffdc8fffedc7;
assign w_fix[58]='h00096afff6f9fffdc2fffdc70001cc;
assign w_fix[59]='hfffe1a000188000338fffe94fffa9c;
assign w_fix[60]='hfffee3fff3c30006ac0011d1fffe8d;
assign w_fix[61]='hfffb4e000544fff816fff9560000d2;
assign w_fix[62]='hfffa450004ba000027fff203000666;
assign w_fix[63]='h00019500004dffffa6001791fffc7e;
assign w_fix[64]='hfffe570010760000fcffff96ffffd0;
assign w_fix[65]='hfff98b0009fb000168001234000058;
assign w_fix[66]='h00008f000d00fffd3a0020b1fffbdc;
assign w_fix[67]='h0002eefffd3c00040ffffaf4ffffb8;
assign w_fix[68]='h0007fb000bca000323fffb6ffffe07;
assign w_fix[69]='hffff63000374000d0cfff5c6000120;
assign w_fix[70]='hffff3dfffe8700007bfffc32000159;
assign w_fix[71]='h0000f1fff7ca0010ee0008d50001ca;
assign w_fix[72]='hfffe7efffb230005d5fff07c0000dc;
assign w_fix[73]='h0000fb000c92000a6cfff7ba000339;
assign w_fix[74]='hfffeb600004cffff25fffee50000f4;
assign w_fix[75]='h000569fffb24000215ffea0a000676;
assign w_fix[76]='hfffc4ffffac2000615ffea13fffe0d;
assign w_fix[77]='hffff67000473fffa510005230001cd;
assign w_fix[78]='hfffd22fffeaffffd9ffff2940003c1;
assign w_fix[79]='h00008e000659fffb16ffee9e0001bb;
assign w_fix[80]='hfffeef000226000ec00007a800027d;
assign w_fix[81]='hfff5ebffff3800042900103c0000b9;
assign w_fix[82]='h000098fffd76ffef3d000bfdfffb4a;
assign w_fix[83]='h0001960003af0003fb0008c1000197;
assign w_fix[84]='h00010effe8910000fc000c2cfffdd3;
assign w_fix[85]='h000159fff27a00067100146a000153;
assign w_fix[86]='hfffffcfff7b000045dffe5c2000011;
assign w_fix[87]='h000097000aa5ffef8fffed47ffffe0;
assign w_fix[88]='h00003b0001da00037e000183000062;
assign w_fix[89]='h0002cdfffc9bffff280000470000c7;
assign w_fix[90]='h000a00000af600014bffdb9d002d89;
assign w_fix[91]='hffffcf0009c90001f7fff645fff7a1;
assign w_fix[92]='h00022c0010f20009c2000c12000bba;
assign w_fix[93]='h00179c00014bfff861ffeb44fffdc0;
assign w_fix[94]='h0000150006c3fffd82fff57afff03b;
assign w_fix[95]='h000aa70009df00276afffea90017a1;
assign w_fix[96]='h0007f8000b160021be0003b2001f60;
assign w_fix[97]='hffff8dffef1f0003c800005600000b;
assign w_fix[98]='hfffe72ffe5c4001546fff6530007fa;
assign w_fix[99]='hfffa700007cdfff84900070cfffb00;
assign w_fix[100]='hfffdf60002edfff9a1fffc90fff85c;
assign w_fix[101]='h0006fa000863001000fff67a000825;
assign w_fix[102]='hfffd32000b88fff6530000f8fff5ac;
assign w_fix[103]='hfff8a7ffec2bfff38e000c26ffde4b;
assign w_fix[104]='h0002460002180000df000147000891;
assign w_fix[105]='hffffd1fff5cbffdf3c000c0effe6bb;
assign w_fix[106]='h0002c6001687ffe7d00004bffff261;
assign w_fix[107]='hfffedc000ddcfffac0fffc0c0011aa;
assign w_fix[108]='h00031500013afff23b000d55ffed1b;
assign w_fix[109]='hffff9afff95cffe97a0006cbffedad;
assign w_fix[110]='hfffe2efffce5000c0ffff80b0019d6;
assign w_fix[111]='hfffc2900201e000289fff8a4000b7f;
assign w_fix[112]='h00131a00130a0031f4fff4c7002bb0;
assign w_fix[113]='h0001990006c600008300095afffbff;
assign w_fix[114]='h0000a6fffa20000628ffc8cc000e60;
assign w_fix[115]='hfffcc9fff8bf000367000cde001429;
assign w_fix[116]='hfff313000850ffed84000badfff38b;
assign w_fix[117]='hfff734fff8a7ffe19f00055effe153;
assign w_fix[118]='h00031900098afff9c1fffecdfffc74;
assign w_fix[119]='h0001fefff5020003440002ac00032a;
assign w_fix[120]='h00096fffe3cc00341ffffc3dfffb76;
assign w_fix[121]='hfff8effff46500037b000e5efffdf8;
assign w_fix[122]='hfff534fff9bb00060300262affeb0c;
assign w_fix[123]='h000f7b000d17fff008000403fff333;
assign w_fix[124]='h000021fff66a00062a00090b000fc5;
assign w_fix[125]='h0002f90018dc002dc7fffa4ffff82f;
assign w_fix[126]='hfff3d300150700279400009b000235;
assign w_fix[127]='h0003710004840002cbfff5d500089c;
assign w_fix[128]='h000388000aa7000c17ffead5000086;
assign w_fix[129]='hfff4bd0002760003b0001407ffffd5;
assign w_fix[130]='hfffd3cfffa08fffde40006e7000092;
assign w_fix[131]='h000d5400086dfff9f4fffdbcfff155;
assign w_fix[132]='hfffc2dfffc86fffe5f0007e1ffff14;
assign w_fix[133]='h0003d9000afcffe45c0001f4fffea6;
assign w_fix[134]='hfffc46ffff14000377000378fffbe4;
assign w_fix[135]='h000431ffebfcffd37f0001f6000750;
assign w_fix[136]='hfff765000371ffee6efffe41fff69f;
assign w_fix[137]='hfff7be000288001e2a000fcdfff960;
assign w_fix[138]='h0002ceffee81ffefdd0012b5000c1d;
assign w_fix[139]='h000159ffef74ffda810001a500151f;
assign w_fix[140]='h0013b000091b004443ffffdf000c39;
assign w_fix[141]='h000c51fffdd3001a92001d6fffef1d;
assign w_fix[142]='h000c0a000bbd001f0bffe962fffaba;
assign w_fix[143]='hfff225fffff900075e000d8e00094e;
assign w_fix[144]='h00097e000737001fc8fffce1ffe9a1;
assign w_fix[145]='h0001df0015bfffec8dfff147fffd49;
assign w_fix[146]='h000415fff3e7fffb48fff982fffb52;
assign w_fix[147]='h0002520004d5ffcf1800112f0004ef;
assign w_fix[148]='hfffa2f00003c0004e1000faf0006a4;
assign w_fix[149]='hffff6500032bfffa16fffddf00001c;
assign w_fix[150]='hfffc8cfffaf90009d0ffef57fff638;
assign w_fix[151]='h00003dfff9cefff73e0006ebfff25d;
assign w_fix[152]='hfffd080001a100035afff6affff0e0;
assign w_fix[153]='hfffdf2001ee1ffee720005b7000903;
assign w_fix[154]='h00006c000034000b2cfffa5dffed75;
assign w_fix[155]='hfffe79000e9200084bfffd5700081b;
assign w_fix[156]='hfffc41000a380009080015f00003b6;
assign w_fix[157]='h00014d000139ffffc400001e0004fb;
assign w_fix[158]='hffffae000112ffd3df000a86fffa73;
assign w_fix[159]='h0001550008bd0003280001ebfffed9;
assign w_fix[160]='h000077000037000330fffa59fffd3f;
assign w_fix[161]='hfffd5e000ccd0007e1000d14fffefb;
assign w_fix[162]='h00016900049d000be2fffb83fffac2;
assign w_fix[163]='h0006ae0001b5000c360005ee0005bf;
assign w_fix[164]='hffff7ffffec3fffad50003890002d4;
assign w_fix[165]='h0002d8fff8f1fff740fffc4dfff876;
assign w_fix[166]='h00026c000fc10019b0fff06a00061f;
assign w_fix[167]='hfffdc300072cfffedb000209001270;
assign w_fix[168]='h00012b00016ffff8010001fbfff8f7;
assign w_fix[169]='hffff49fffb34fffe60000867fffea5;
assign w_fix[170]='h0002b1000c650013550001baffedef;
assign w_fix[171]='hfffdc1000c1a001632fffc79ffec90;
assign w_fix[172]='hfffaebfffe1a000186001133fffcd6;
assign w_fix[173]='h0000ec00064bfff6c4fffc6b000228;
assign w_fix[174]='hffff1e000276ffec7bfff896ffffba;
assign w_fix[175]='hffff5f000aa2000523ffffc4001149;
assign w_fix[176]='h00005a00006b002204fffb840004e4;
assign w_fix[177]='h00021c000381fff46afffa8c000557;
assign w_fix[178]='h0001660002ccfffa6f000056000462;
assign w_fix[179]='h0001bcffffbaffedfc00045e000875;

endmodule