module createAandB_tanh #(
parameter aDW = 18,
parameter bDW = 18,
parameter numOfDots = 549, //�����зֵ�ĸ������������Ҷ˵�
parameter MW = 10
)(
input wire en,
input wire rst_n,
input wire [MW : 0] i,
output reg [(aDW - 1) : 0] a,
output reg [(bDW - 1) : 0] b
);

wire EN;

wire [(aDW - 1) : 0] aList [(numOfDots - 1) : 0];
wire [(bDW - 1) : 0] bList [(numOfDots - 1) : 0];

// assign aList[0] = 16'h0000; 
// assign aList[1] = 16'h0005; 
// assign aList[2] = 16'h004b; 
// assign aList[3] = 16'h00cd; 
// assign aList[4] = 16'h01a3; 
// assign aList[5] = 16'h02b0; 
// assign aList[6] = 16'h0466; 
// assign aList[7] = 16'h064d; 
// assign aList[8] = 16'h0809; 
// assign aList[9] = 16'h0a39; 
// assign aList[10] = 16'h0cf9; 
// assign aList[11] = 16'h106a; 
// assign aList[12] = 16'h14af; 
// assign aList[13] = 16'h19ee; 
// assign aList[14] = 16'h1e8e; 
// assign aList[15] = 16'h220b; 
// assign aList[16] = 16'h25da; 
// assign aList[17] = 16'h29fc; 
// assign aList[18] = 16'h2e74; 
// assign aList[19] = 16'h3340; 
// assign aList[20] = 16'h385e; 
// assign aList[21] = 16'h3dc8; 
// assign aList[22] = 16'h4375; 
// assign aList[23] = 16'h495b; 
// assign aList[24] = 16'h4f69; 
// assign aList[25] = 16'h558e; 
// assign aList[26] = 16'h5bb0; 
// assign aList[27] = 16'h61b7; 
// assign aList[28] = 16'h6785; 
// assign aList[29] = 16'h6cfb; 
// assign aList[30] = 16'h71f7; 
// assign aList[31] = 16'h765b; 
// assign aList[32] = 16'h7b76; 
// assign aList[33] = 16'h7f56; 
// assign aList[34] = 16'h7f56; 
// assign aList[35] = 16'h7b76; 
// assign aList[36] = 16'h765b; 
// assign aList[37] = 16'h71f7; 
// assign aList[38] = 16'h6cfb; 
// assign aList[39] = 16'h6785; 
// assign aList[40] = 16'h61b7; 
// assign aList[41] = 16'h5bb0; 
// assign aList[42] = 16'h558e; 
// assign aList[43] = 16'h4f69; 
// assign aList[44] = 16'h495b; 
// assign aList[45] = 16'h4375; 
// assign aList[46] = 16'h3dc8; 
// assign aList[47] = 16'h385e; 
// assign aList[48] = 16'h3340; 
// assign aList[49] = 16'h2e74; 
// assign aList[50] = 16'h29fc; 
// assign aList[51] = 16'h25da; 
// assign aList[52] = 16'h220b; 
// assign aList[53] = 16'h1e8e; 
// assign aList[54] = 16'h19ee; 
// assign aList[55] = 16'h14af; 
// assign aList[56] = 16'h106a; 
// assign aList[57] = 16'h0cf9; 
// assign aList[58] = 16'h0a39; 
// assign aList[59] = 16'h0809; 
// assign aList[60] = 16'h064d; 
// assign aList[61] = 16'h0466; 
// assign aList[62] = 16'h02b0; 
// assign aList[63] = 16'h01a3; 
// assign aList[64] = 16'h00cd; 
// assign aList[65] = 16'h004b; 
// assign aList[66] = 16'h0005; 

// assign bList[0] = 16'h0000;
// assign bList[1] = 16'h802c; 
// assign bList[2] = 16'h8144; 
// assign bList[3] = 16'h8308; 
// assign bList[4] = 16'h858a; 
// assign bList[5] = 16'h886d; 
// assign bList[6] = 16'h8cb5; 
// assign bList[7] = 16'h90fd; 
// assign bList[8] = 16'h94ac; 
// assign bList[9] = 16'h990c; 
// assign bList[10] = 16'h9e35; 
// assign bList[11] = 16'ha43a; 
// assign bList[12] = 16'hab2a; 
// assign bList[13] = 16'hb309; 
// assign bList[14] = 16'hb966; 
// assign bList[15] = 16'hbdf9; 
// assign bList[16] = 16'hc2bc; 
// assign bList[17] = 16'hc7a5; 
// assign bList[18] = 16'hccab; 
// assign bList[19] = 16'hd1c4; 
// assign bList[20] = 16'hd6e2; 
// assign bList[21] = 16'hdbf5; 
// assign bList[22] = 16'he0ed; 
// assign bList[23] = 16'he5b8; 
// assign bList[24] = 16'hea43; 
// assign bList[25] = 16'hee7b; 
// assign bList[26] = 16'hf251; 
// assign bList[27] = 16'hf5b5; 
// assign bList[28] = 16'hf89c; 
// assign bList[29] = 16'hfaff; 
// assign bList[30] = 16'hfcde; 
// assign bList[31] = 16'hfe3d; 
// assign bList[32] = 16'hff84; 
// assign bList[33] = 16'h0000; 
// assign bList[34] = 16'h0000; 
// assign bList[35] = 16'h007c; 
// assign bList[36] = 16'h01c3; 
// assign bList[37] = 16'h0322; 
// assign bList[38] = 16'h0501; 
// assign bList[39] = 16'h0764; 
// assign bList[40] = 16'h0a4b; 
// assign bList[41] = 16'h0daf; 
// assign bList[42] = 16'h1185; 
// assign bList[43] = 16'h15bd; 
// assign bList[44] = 16'h1a48; 
// assign bList[45] = 16'h1f13; 
// assign bList[46] = 16'h240b; 
// assign bList[47] = 16'h291e; 
// assign bList[48] = 16'h2e3c; 
// assign bList[49] = 16'h3355; 
// assign bList[50] = 16'h385b; 
// assign bList[51] = 16'h3d44; 
// assign bList[52] = 16'h4207; 
// assign bList[53] = 16'h469a; 
// assign bList[54] = 16'h4cf7; 
// assign bList[55] = 16'h54d6; 
// assign bList[56] = 16'h5bc6; 
// assign bList[57] = 16'h61cb; 
// assign bList[58] = 16'h66f4; 
// assign bList[59] = 16'h6b54; 
// assign bList[60] = 16'h6f03; 
// assign bList[61] = 16'h734b; 
// assign bList[62] = 16'h7793; 
// assign bList[63] = 16'h7a76; 
// assign bList[64] = 16'h7cf8; 
// assign bList[65] = 16'h7ebc; 
// assign bList[66] = 16'h7fd4; 

assign aList[0] = 18'h00000; 
assign aList[1] = 18'h00001; 
assign aList[2] = 18'h00006; 
assign aList[3] = 18'h0000f; 
assign aList[4] = 18'h0001f; 
assign aList[5] = 18'h00033; 
assign aList[6] = 18'h00054; 
assign aList[7] = 18'h00079; 
assign aList[8] = 18'h0009c; 
assign aList[9] = 18'h000c8; 
assign aList[10] = 18'h00100; 
assign aList[11] = 18'h00149; 
assign aList[12] = 18'h0018c; 
assign aList[13] = 18'h001c1; 
assign aList[14] = 18'h001fc; 
assign aList[15] = 18'h00240; 
assign aList[16] = 18'h0028c; 
assign aList[17] = 18'h002e3; 
assign aList[18] = 18'h00345; 
assign aList[19] = 18'h003b4; 
assign aList[20] = 18'h00432; 
assign aList[21] = 18'h004c0; 
assign aList[22] = 18'h00536; 
assign aList[23] = 18'h0058c; 
assign aList[24] = 18'h005e7; 
assign aList[25] = 18'h00648; 
assign aList[26] = 18'h006af; 
assign aList[27] = 18'h0071c; 
assign aList[28] = 18'h00791; 
assign aList[29] = 18'h0080d; 
assign aList[30] = 18'h00890; 
assign aList[31] = 18'h0091d; 
assign aList[32] = 18'h009b2; 
assign aList[33] = 18'h00a50; 
assign aList[34] = 18'h00af8; 
assign aList[35] = 18'h00bac; 
assign aList[36] = 18'h00c6a; 
assign aList[37] = 18'h00d34; 
assign aList[38] = 18'h00e0b; 
assign aList[39] = 18'h00ef0; 
assign aList[40] = 18'h00fe2; 
assign aList[41] = 18'h010e4; 
assign aList[42] = 18'h011f6; 
assign aList[43] = 18'h01319; 
assign aList[44] = 18'h0144e; 
assign aList[45] = 18'h01542; 
assign aList[46] = 18'h015eb; 
assign aList[47] = 18'h01699; 
assign aList[48] = 18'h0174c; 
assign aList[49] = 18'h01805; 
assign aList[50] = 18'h018c4; 
assign aList[51] = 18'h01988; 
assign aList[52] = 18'h01a52; 
assign aList[53] = 18'h01b22; 
assign aList[54] = 18'h01bf8; 
assign aList[55] = 18'h01cd5; 
assign aList[56] = 18'h01db9; 
assign aList[57] = 18'h01ea3; 
assign aList[58] = 18'h01f94; 
assign aList[59] = 18'h0208c; 
assign aList[60] = 18'h0218c; 
assign aList[61] = 18'h02293; 
assign aList[62] = 18'h023a2; 
assign aList[63] = 18'h024b9; 
assign aList[64] = 18'h025d8; 
assign aList[65] = 18'h02700; 
assign aList[66] = 18'h02830; 
assign aList[67] = 18'h02969; 
assign aList[68] = 18'h02aac; 
assign aList[69] = 18'h02bf7; 
assign aList[70] = 18'h02d4c; 
assign aList[71] = 18'h02eab; 
assign aList[72] = 18'h03014; 
assign aList[73] = 18'h03187; 
assign aList[74] = 18'h03305; 
assign aList[75] = 18'h0348e; 
assign aList[76] = 18'h03622; 
assign aList[77] = 18'h037c1; 
assign aList[78] = 18'h0396c; 
assign aList[79] = 18'h03b23; 
assign aList[80] = 18'h03ce6; 
assign aList[81] = 18'h03eb6; 
assign aList[82] = 18'h04092; 
assign aList[83] = 18'h0427c; 
assign aList[84] = 18'h04472; 
assign aList[85] = 18'h04677; 
assign aList[86] = 18'h0488a; 
assign aList[87] = 18'h04aaa; 
assign aList[88] = 18'h04cda; 
assign aList[89] = 18'h04f18; 
assign aList[90] = 18'h05166; 
assign aList[91] = 18'h053c2; 
assign aList[92] = 18'h0562f; 
assign aList[93] = 18'h058ac; 
assign aList[94] = 18'h05b39; 
assign aList[95] = 18'h05d2e; 
assign aList[96] = 18'h05e81; 
assign aList[97] = 18'h05fd8; 
assign aList[98] = 18'h06134; 
assign aList[99] = 18'h06294; 
assign aList[100] = 18'h063f9; 
assign aList[101] = 18'h06562; 
assign aList[102] = 18'h066cf; 
assign aList[103] = 18'h06841; 
assign aList[104] = 18'h069b8; 
assign aList[105] = 18'h06b33; 
assign aList[106] = 18'h06cb2; 
assign aList[107] = 18'h06e36; 
assign aList[108] = 18'h06fbf; 
assign aList[109] = 18'h0714d; 
assign aList[110] = 18'h072df; 
assign aList[111] = 18'h07476; 
assign aList[112] = 18'h07612; 
assign aList[113] = 18'h077b3; 
assign aList[114] = 18'h07958; 
assign aList[115] = 18'h07b03; 
assign aList[116] = 18'h07cb2; 
assign aList[117] = 18'h07e66; 
assign aList[118] = 18'h08020; 
assign aList[119] = 18'h081de; 
assign aList[120] = 18'h083a1; 
assign aList[121] = 18'h08569; 
assign aList[122] = 18'h08737; 
assign aList[123] = 18'h08909; 
assign aList[124] = 18'h08ae1; 
assign aList[125] = 18'h08cbe; 
assign aList[126] = 18'h08ea0; 
assign aList[127] = 18'h09087; 
assign aList[128] = 18'h09273; 
assign aList[129] = 18'h09465; 
assign aList[130] = 18'h0965c; 
assign aList[131] = 18'h09858; 
assign aList[132] = 18'h09a59; 
assign aList[133] = 18'h09c60; 
assign aList[134] = 18'h09e6c; 
assign aList[135] = 18'h0a07d; 
assign aList[136] = 18'h0a294; 
assign aList[137] = 18'h0a4b0; 
assign aList[138] = 18'h0a6d1; 
assign aList[139] = 18'h0a8f7; 
assign aList[140] = 18'h0ab23; 
assign aList[141] = 18'h0ad54; 
assign aList[142] = 18'h0af8b; 
assign aList[143] = 18'h0b1c7; 
assign aList[144] = 18'h0b408; 
assign aList[145] = 18'h0b64f; 
assign aList[146] = 18'h0b89a; 
assign aList[147] = 18'h0baeb; 
assign aList[148] = 18'h0bd42; 
assign aList[149] = 18'h0bf9e; 
assign aList[150] = 18'h0c1fe; 
assign aList[151] = 18'h0c465; 
assign aList[152] = 18'h0c6d0; 
assign aList[153] = 18'h0c941; 
assign aList[154] = 18'h0cbb6; 
assign aList[155] = 18'h0ce31; 
assign aList[156] = 18'h0d0b1; 
assign aList[157] = 18'h0d336; 
assign aList[158] = 18'h0d5c0; 
assign aList[159] = 18'h0d84f; 
assign aList[160] = 18'h0dae3; 
assign aList[161] = 18'h0dd7c; 
assign aList[162] = 18'h0e01a; 
assign aList[163] = 18'h0e2bc; 
assign aList[164] = 18'h0e564; 
assign aList[165] = 18'h0e810; 
assign aList[166] = 18'h0eac1; 
assign aList[167] = 18'h0ed76; 
assign aList[168] = 18'h0f030; 
assign aList[169] = 18'h0f2ee; 
assign aList[170] = 18'h0f5b0; 
assign aList[171] = 18'h0f877; 
assign aList[172] = 18'h0fb42; 
assign aList[173] = 18'h0fe12; 
assign aList[174] = 18'h100e5; 
assign aList[175] = 18'h103bc; 
assign aList[176] = 18'h10698; 
assign aList[177] = 18'h10976; 
assign aList[178] = 18'h10c59; 
assign aList[179] = 18'h10f3f; 
assign aList[180] = 18'h11229; 
assign aList[181] = 18'h11516; 
assign aList[182] = 18'h11807; 
assign aList[183] = 18'h11afa; 
assign aList[184] = 18'h11df1; 
assign aList[185] = 18'h120ea; 
assign aList[186] = 18'h123e6; 
assign aList[187] = 18'h126e5; 
assign aList[188] = 18'h129e6; 
assign aList[189] = 18'h12cea; 
assign aList[190] = 18'h12ff0; 
assign aList[191] = 18'h132f8; 
assign aList[192] = 18'h13602; 
assign aList[193] = 18'h1390e; 
assign aList[194] = 18'h13c1b; 
assign aList[195] = 18'h13f2a; 
assign aList[196] = 18'h1423a; 
assign aList[197] = 18'h1454b; 
assign aList[198] = 18'h1485d; 
assign aList[199] = 18'h14b70; 
assign aList[200] = 18'h14e84; 
assign aList[201] = 18'h15198; 
assign aList[202] = 18'h154ac; 
assign aList[203] = 18'h157c0; 
assign aList[204] = 18'h15ad4; 
assign aList[205] = 18'h15de8; 
assign aList[206] = 18'h160fb; 
assign aList[207] = 18'h1640e; 
assign aList[208] = 18'h1671f; 
assign aList[209] = 18'h16a30; 
assign aList[210] = 18'h16d3f; 
assign aList[211] = 18'h1704c; 
assign aList[212] = 18'h17357; 
assign aList[213] = 18'h17661; 
assign aList[214] = 18'h17968; 
assign aList[215] = 18'h17c6d; 
assign aList[216] = 18'h17f6f; 
assign aList[217] = 18'h1826e; 
assign aList[218] = 18'h1856a; 
assign aList[219] = 18'h18862; 
assign aList[220] = 18'h18b57; 
assign aList[221] = 18'h18e48; 
assign aList[222] = 18'h19134; 
assign aList[223] = 18'h1941d; 
assign aList[224] = 18'h19700; 
assign aList[225] = 18'h199df; 
assign aList[226] = 18'h19cb9; 
assign aList[227] = 18'h19f8d; 
assign aList[228] = 18'h1a25b; 
assign aList[229] = 18'h1a524; 
assign aList[230] = 18'h1a7e7; 
assign aList[231] = 18'h1aaa3; 
assign aList[232] = 18'h1ad58; 
assign aList[233] = 18'h1b007; 
assign aList[234] = 18'h1b2ae; 
assign aList[235] = 18'h1b54e; 
assign aList[236] = 18'h1b7e6; 
assign aList[237] = 18'h1ba76; 
assign aList[238] = 18'h1bcfe; 
assign aList[239] = 18'h1bf7e; 
assign aList[240] = 18'h1c1f5; 
assign aList[241] = 18'h1c463; 
assign aList[242] = 18'h1c6c8; 
assign aList[243] = 18'h1c923; 
assign aList[244] = 18'h1cb75; 
assign aList[245] = 18'h1cdbd; 
assign aList[246] = 18'h1cffa; 
assign aList[247] = 18'h1d22d; 
assign aList[248] = 18'h1d456; 
assign aList[249] = 18'h1d673; 
assign aList[250] = 18'h1d886; 
assign aList[251] = 18'h1da8d; 
assign aList[252] = 18'h1dc88; 
assign aList[253] = 18'h1de78; 
assign aList[254] = 18'h1e05c; 
assign aList[255] = 18'h1e233; 
assign aList[256] = 18'h1e3fe; 
assign aList[257] = 18'h1e5bd; 
assign aList[258] = 18'h1e76e; 
assign aList[259] = 18'h1e913; 
assign aList[260] = 18'h1eaaa; 
assign aList[261] = 18'h1ec34; 
assign aList[262] = 18'h1edb0; 
assign aList[263] = 18'h1ef1f; 
assign aList[264] = 18'h1f07f; 
assign aList[265] = 18'h1f274; 
assign aList[266] = 18'h1f4df; 
assign aList[267] = 18'h1f710; 
assign aList[268] = 18'h1f906; 
assign aList[269] = 18'h1fabf; 
assign aList[270] = 18'h1fc3a; 
assign aList[271] = 18'h1fd78; 
assign aList[272] = 18'h1fe76; 
assign aList[273] = 18'h1ff36; 
assign aList[274] = 18'h1ffd5; 
assign aList[275] = 18'h1ffd5; 
assign aList[276] = 18'h1ff36; 
assign aList[277] = 18'h1fe76; 
assign aList[278] = 18'h1fd78; 
assign aList[279] = 18'h1fc3a; 
assign aList[280] = 18'h1fabf; 
assign aList[281] = 18'h1f906; 
assign aList[282] = 18'h1f710; 
assign aList[283] = 18'h1f4df; 
assign aList[284] = 18'h1f274; 
assign aList[285] = 18'h1f07f; 
assign aList[286] = 18'h1ef1f; 
assign aList[287] = 18'h1edb0; 
assign aList[288] = 18'h1ec34; 
assign aList[289] = 18'h1eaaa; 
assign aList[290] = 18'h1e913; 
assign aList[291] = 18'h1e76e; 
assign aList[292] = 18'h1e5bd; 
assign aList[293] = 18'h1e3fe; 
assign aList[294] = 18'h1e233; 
assign aList[295] = 18'h1e05c; 
assign aList[296] = 18'h1de78; 
assign aList[297] = 18'h1dc88; 
assign aList[298] = 18'h1da8d; 
assign aList[299] = 18'h1d886; 
assign aList[300] = 18'h1d673; 
assign aList[301] = 18'h1d456; 
assign aList[302] = 18'h1d22d; 
assign aList[303] = 18'h1cffa; 
assign aList[304] = 18'h1cdbd; 
assign aList[305] = 18'h1cb75; 
assign aList[306] = 18'h1c923; 
assign aList[307] = 18'h1c6c8; 
assign aList[308] = 18'h1c463; 
assign aList[309] = 18'h1c1f5; 
assign aList[310] = 18'h1bf7e; 
assign aList[311] = 18'h1bcfe; 
assign aList[312] = 18'h1ba76; 
assign aList[313] = 18'h1b7e6; 
assign aList[314] = 18'h1b54e; 
assign aList[315] = 18'h1b2ae; 
assign aList[316] = 18'h1b007; 
assign aList[317] = 18'h1ad58; 
assign aList[318] = 18'h1aaa3; 
assign aList[319] = 18'h1a7e7; 
assign aList[320] = 18'h1a524; 
assign aList[321] = 18'h1a25b; 
assign aList[322] = 18'h19f8d; 
assign aList[323] = 18'h19cb9; 
assign aList[324] = 18'h199df; 
assign aList[325] = 18'h19700; 
assign aList[326] = 18'h1941d; 
assign aList[327] = 18'h19134; 
assign aList[328] = 18'h18e48; 
assign aList[329] = 18'h18b57; 
assign aList[330] = 18'h18862; 
assign aList[331] = 18'h1856a; 
assign aList[332] = 18'h1826e; 
assign aList[333] = 18'h17f6f; 
assign aList[334] = 18'h17c6d; 
assign aList[335] = 18'h17968; 
assign aList[336] = 18'h17661; 
assign aList[337] = 18'h17357; 
assign aList[338] = 18'h1704c; 
assign aList[339] = 18'h16d3f; 
assign aList[340] = 18'h16a30; 
assign aList[341] = 18'h1671f; 
assign aList[342] = 18'h1640e; 
assign aList[343] = 18'h160fb; 
assign aList[344] = 18'h15de8; 
assign aList[345] = 18'h15ad4; 
assign aList[346] = 18'h157c0; 
assign aList[347] = 18'h154ac; 
assign aList[348] = 18'h15198; 
assign aList[349] = 18'h14e84; 
assign aList[350] = 18'h14b70; 
assign aList[351] = 18'h1485d; 
assign aList[352] = 18'h1454b; 
assign aList[353] = 18'h1423a; 
assign aList[354] = 18'h13f2a; 
assign aList[355] = 18'h13c1b; 
assign aList[356] = 18'h1390e; 
assign aList[357] = 18'h13602; 
assign aList[358] = 18'h132f8; 
assign aList[359] = 18'h12ff0; 
assign aList[360] = 18'h12cea; 
assign aList[361] = 18'h129e6; 
assign aList[362] = 18'h126e5; 
assign aList[363] = 18'h123e6; 
assign aList[364] = 18'h120ea; 
assign aList[365] = 18'h11df1; 
assign aList[366] = 18'h11afa; 
assign aList[367] = 18'h11807; 
assign aList[368] = 18'h11516; 
assign aList[369] = 18'h11229; 
assign aList[370] = 18'h10f3f; 
assign aList[371] = 18'h10c59; 
assign aList[372] = 18'h10976; 
assign aList[373] = 18'h10698; 
assign aList[374] = 18'h103bc; 
assign aList[375] = 18'h100e5; 
assign aList[376] = 18'h0fe12; 
assign aList[377] = 18'h0fb42; 
assign aList[378] = 18'h0f877; 
assign aList[379] = 18'h0f5b0; 
assign aList[380] = 18'h0f2ee; 
assign aList[381] = 18'h0f030; 
assign aList[382] = 18'h0ed76; 
assign aList[383] = 18'h0eac1; 
assign aList[384] = 18'h0e810; 
assign aList[385] = 18'h0e564; 
assign aList[386] = 18'h0e2bc; 
assign aList[387] = 18'h0e01a; 
assign aList[388] = 18'h0dd7c; 
assign aList[389] = 18'h0dae3; 
assign aList[390] = 18'h0d84f; 
assign aList[391] = 18'h0d5c0; 
assign aList[392] = 18'h0d336; 
assign aList[393] = 18'h0d0b1; 
assign aList[394] = 18'h0ce31; 
assign aList[395] = 18'h0cbb6; 
assign aList[396] = 18'h0c941; 
assign aList[397] = 18'h0c6d0; 
assign aList[398] = 18'h0c465; 
assign aList[399] = 18'h0c1fe; 
assign aList[400] = 18'h0bf9e; 
assign aList[401] = 18'h0bd42; 
assign aList[402] = 18'h0baeb; 
assign aList[403] = 18'h0b89a; 
assign aList[404] = 18'h0b64f; 
assign aList[405] = 18'h0b408; 
assign aList[406] = 18'h0b1c7; 
assign aList[407] = 18'h0af8b; 
assign aList[408] = 18'h0ad54; 
assign aList[409] = 18'h0ab23; 
assign aList[410] = 18'h0a8f7; 
assign aList[411] = 18'h0a6d1; 
assign aList[412] = 18'h0a4b0; 
assign aList[413] = 18'h0a294; 
assign aList[414] = 18'h0a07d; 
assign aList[415] = 18'h09e6c; 
assign aList[416] = 18'h09c60; 
assign aList[417] = 18'h09a59; 
assign aList[418] = 18'h09858; 
assign aList[419] = 18'h0965c; 
assign aList[420] = 18'h09465; 
assign aList[421] = 18'h09273; 
assign aList[422] = 18'h09087; 
assign aList[423] = 18'h08ea0; 
assign aList[424] = 18'h08cbe; 
assign aList[425] = 18'h08ae1; 
assign aList[426] = 18'h08909; 
assign aList[427] = 18'h08737; 
assign aList[428] = 18'h08569; 
assign aList[429] = 18'h083a1; 
assign aList[430] = 18'h081de; 
assign aList[431] = 18'h08020; 
assign aList[432] = 18'h07e66; 
assign aList[433] = 18'h07cb2; 
assign aList[434] = 18'h07b03; 
assign aList[435] = 18'h07958; 
assign aList[436] = 18'h077b3; 
assign aList[437] = 18'h07612; 
assign aList[438] = 18'h07476; 
assign aList[439] = 18'h072df; 
assign aList[440] = 18'h0714d; 
assign aList[441] = 18'h06fbf; 
assign aList[442] = 18'h06e36; 
assign aList[443] = 18'h06cb2; 
assign aList[444] = 18'h06b33; 
assign aList[445] = 18'h069b8; 
assign aList[446] = 18'h06841; 
assign aList[447] = 18'h066cf; 
assign aList[448] = 18'h06562; 
assign aList[449] = 18'h063f9; 
assign aList[450] = 18'h06294; 
assign aList[451] = 18'h06134; 
assign aList[452] = 18'h05fd8; 
assign aList[453] = 18'h05e81; 
assign aList[454] = 18'h05d2e; 
assign aList[455] = 18'h05b39; 
assign aList[456] = 18'h058ac; 
assign aList[457] = 18'h0562f; 
assign aList[458] = 18'h053c2; 
assign aList[459] = 18'h05166; 
assign aList[460] = 18'h04f18; 
assign aList[461] = 18'h04cda; 
assign aList[462] = 18'h04aaa; 
assign aList[463] = 18'h0488a; 
assign aList[464] = 18'h04677; 
assign aList[465] = 18'h04472; 
assign aList[466] = 18'h0427c; 
assign aList[467] = 18'h04092; 
assign aList[468] = 18'h03eb6; 
assign aList[469] = 18'h03ce6; 
assign aList[470] = 18'h03b23; 
assign aList[471] = 18'h0396c; 
assign aList[472] = 18'h037c1; 
assign aList[473] = 18'h03622; 
assign aList[474] = 18'h0348e; 
assign aList[475] = 18'h03305; 
assign aList[476] = 18'h03187; 
assign aList[477] = 18'h03014; 
assign aList[478] = 18'h02eab; 
assign aList[479] = 18'h02d4c; 
assign aList[480] = 18'h02bf7; 
assign aList[481] = 18'h02aac; 
assign aList[482] = 18'h02969; 
assign aList[483] = 18'h02830; 
assign aList[484] = 18'h02700; 
assign aList[485] = 18'h025d8; 
assign aList[486] = 18'h024b9; 
assign aList[487] = 18'h023a2; 
assign aList[488] = 18'h02293; 
assign aList[489] = 18'h0218c; 
assign aList[490] = 18'h0208c; 
assign aList[491] = 18'h01f94; 
assign aList[492] = 18'h01ea3; 
assign aList[493] = 18'h01db9; 
assign aList[494] = 18'h01cd5; 
assign aList[495] = 18'h01bf8; 
assign aList[496] = 18'h01b22; 
assign aList[497] = 18'h01a52; 
assign aList[498] = 18'h01988; 
assign aList[499] = 18'h018c4; 
assign aList[500] = 18'h01805; 
assign aList[501] = 18'h0174c; 
assign aList[502] = 18'h01699; 
assign aList[503] = 18'h015eb; 
assign aList[504] = 18'h01542; 
assign aList[505] = 18'h0144e; 
assign aList[506] = 18'h01319; 
assign aList[507] = 18'h011f6; 
assign aList[508] = 18'h010e4; 
assign aList[509] = 18'h00fe2; 
assign aList[510] = 18'h00ef0; 
assign aList[511] = 18'h00e0b; 
assign aList[512] = 18'h00d34; 
assign aList[513] = 18'h00c6a; 
assign aList[514] = 18'h00bac; 
assign aList[515] = 18'h00af8; 
assign aList[516] = 18'h00a50; 
assign aList[517] = 18'h009b2; 
assign aList[518] = 18'h0091d; 
assign aList[519] = 18'h00890; 
assign aList[520] = 18'h0080d; 
assign aList[521] = 18'h00791; 
assign aList[522] = 18'h0071c; 
assign aList[523] = 18'h006af; 
assign aList[524] = 18'h00648; 
assign aList[525] = 18'h005e7; 
assign aList[526] = 18'h0058c; 
assign aList[527] = 18'h00536; 
assign aList[528] = 18'h004c0; 
assign aList[529] = 18'h00432; 
assign aList[530] = 18'h003b4; 
assign aList[531] = 18'h00345; 
assign aList[532] = 18'h002e3; 
assign aList[533] = 18'h0028c; 
assign aList[534] = 18'h00240; 
assign aList[535] = 18'h001fc; 
assign aList[536] = 18'h001c1; 
assign aList[537] = 18'h0018c; 
assign aList[538] = 18'h00149; 
assign aList[539] = 18'h00100; 
assign aList[540] = 18'h000c8; 
assign aList[541] = 18'h0009c; 
assign aList[542] = 18'h00079; 
assign aList[543] = 18'h00054; 
assign aList[544] = 18'h00033; 
assign aList[545] = 18'h0001f; 
assign aList[546] = 18'h0000f; 
assign aList[547] = 18'h00006; 
assign aList[548] = 18'h00001; 

assign bList[0] = 18'h00000; 
assign bList[1] = 18'h20006; 
assign bList[2] = 18'h20023; 
assign bList[3] = 18'h20057; 
assign bList[4] = 18'h200a6; 
assign bList[5] = 18'h20105; 
assign bList[6] = 18'h2019a; 
assign bList[7] = 18'h20238; 
assign bList[8] = 18'h202c6; 
assign bList[9] = 18'h20377; 
assign bList[10] = 18'h20452; 
assign bList[11] = 18'h20563; 
assign bList[12] = 18'h20656; 
assign bList[13] = 18'h20711; 
assign bList[14] = 18'h207e2; 
assign bList[15] = 18'h208ca; 
assign bList[16] = 18'h209cc; 
assign bList[17] = 18'h20aeb; 
assign bList[18] = 18'h20c2a; 
assign bList[19] = 18'h20d8b; 
assign bList[20] = 18'h20f14; 
assign bList[21] = 18'h210c8; 
assign bList[22] = 18'h2122b; 
assign bList[23] = 18'h21329; 
assign bList[24] = 18'h21434; 
assign bList[25] = 18'h2154e; 
assign bList[26] = 18'h21676; 
assign bList[27] = 18'h217ad; 
assign bList[28] = 18'h218f5; 
assign bList[29] = 18'h21a4e; 
assign bList[30] = 18'h21bb8; 
assign bList[31] = 18'h21d35; 
assign bList[32] = 18'h21ec6; 
assign bList[33] = 18'h2206b; 
assign bList[34] = 18'h22225; 
assign bList[35] = 18'h223f5; 
assign bList[36] = 18'h225dd; 
assign bList[37] = 18'h227dd; 
assign bList[38] = 18'h229f6; 
assign bList[39] = 18'h22c2a; 
assign bList[40] = 18'h22e7a; 
assign bList[41] = 18'h230e7; 
assign bList[42] = 18'h23371; 
assign bList[43] = 18'h2361b; 
assign bList[44] = 18'h238e6; 
assign bList[45] = 18'h23b12; 
assign bList[46] = 18'h23c91; 
assign bList[47] = 18'h23e18; 
assign bList[48] = 18'h23fa9; 
assign bList[49] = 18'h24143; 
assign bList[50] = 18'h242e7; 
assign bList[51] = 18'h24494; 
assign bList[52] = 18'h2464b; 
assign bList[53] = 18'h2480c; 
assign bList[54] = 18'h249d6; 
assign bList[55] = 18'h24bac; 
assign bList[56] = 18'h24d8b; 
assign bList[57] = 18'h24f76; 
assign bList[58] = 18'h2516b; 
assign bList[59] = 18'h2536b; 
assign bList[60] = 18'h25576; 
assign bList[61] = 18'h2578d; 
assign bList[62] = 18'h259af; 
assign bList[63] = 18'h25bdd; 
assign bList[64] = 18'h25e17; 
assign bList[65] = 18'h2605d; 
assign bList[66] = 18'h262af; 
assign bList[67] = 18'h2650e; 
assign bList[68] = 18'h26779; 
assign bList[69] = 18'h269f1; 
assign bList[70] = 18'h26c76; 
assign bList[71] = 18'h26f08; 
assign bList[72] = 18'h271a7; 
assign bList[73] = 18'h27454; 
assign bList[74] = 18'h2770e; 
assign bList[75] = 18'h279d6; 
assign bList[76] = 18'h27cac; 
assign bList[77] = 18'h27f90; 
assign bList[78] = 18'h28281; 
assign bList[79] = 18'h28581; 
assign bList[80] = 18'h28890; 
assign bList[81] = 18'h28bac; 
assign bList[82] = 18'h28ed8; 
assign bList[83] = 18'h29212; 
assign bList[84] = 18'h2955b; 
assign bList[85] = 18'h298b2; 
assign bList[86] = 18'h29c19; 
assign bList[87] = 18'h29f8e; 
assign bList[88] = 18'h2a312; 
assign bList[89] = 18'h2a6a5; 
assign bList[90] = 18'h2aa48; 
assign bList[91] = 18'h2adf9; 
assign bList[92] = 18'h2b1b9; 
assign bList[93] = 18'h2b588; 
assign bList[94] = 18'h2b966; 
assign bList[95] = 18'h2bc55; 
assign bList[96] = 18'h2be4f; 
assign bList[97] = 18'h2c04d; 
assign bList[98] = 18'h2c24f; 
assign bList[99] = 18'h2c454; 
assign bList[100] = 18'h2c65d; 
assign bList[101] = 18'h2c869; 
assign bList[102] = 18'h2ca79; 
assign bList[103] = 18'h2cc8d; 
assign bList[104] = 18'h2cea4; 
assign bList[105] = 18'h2d0bf; 
assign bList[106] = 18'h2d2de; 
assign bList[107] = 18'h2d500; 
assign bList[108] = 18'h2d725; 
assign bList[109] = 18'h2d94e; 
assign bList[110] = 18'h2db7a; 
assign bList[111] = 18'h2ddaa; 
assign bList[112] = 18'h2dfdd; 
assign bList[113] = 18'h2e213; 
assign bList[114] = 18'h2e44d; 
assign bList[115] = 18'h2e68a; 
assign bList[116] = 18'h2e8ca; 
assign bList[117] = 18'h2eb0e; 
assign bList[118] = 18'h2ed54; 
assign bList[119] = 18'h2ef9e; 
assign bList[120] = 18'h2f1eb; 
assign bList[121] = 18'h2f43b; 
assign bList[122] = 18'h2f68d; 
assign bList[123] = 18'h2f8e3; 
assign bList[124] = 18'h2fb3c; 
assign bList[125] = 18'h2fd97; 
assign bList[126] = 18'h2fff6; 
assign bList[127] = 18'h30256; 
assign bList[128] = 18'h304ba; 
assign bList[129] = 18'h30720; 
assign bList[130] = 18'h30989; 
assign bList[131] = 18'h30bf4; 
assign bList[132] = 18'h30e62; 
assign bList[133] = 18'h310d2; 
assign bList[134] = 18'h31344; 
assign bList[135] = 18'h315b9; 
assign bList[136] = 18'h3182f; 
assign bList[137] = 18'h31aa8; 
assign bList[138] = 18'h31d23; 
assign bList[139] = 18'h31f9f; 
assign bList[140] = 18'h3221e; 
assign bList[141] = 18'h3249e; 
assign bList[142] = 18'h32720; 
assign bList[143] = 18'h329a3; 
assign bList[144] = 18'h32c28; 
assign bList[145] = 18'h32eae; 
assign bList[146] = 18'h33136; 
assign bList[147] = 18'h333be; 
assign bList[148] = 18'h33648; 
assign bList[149] = 18'h338d3; 
assign bList[150] = 18'h33b5f; 
assign bList[151] = 18'h33deb; 
assign bList[152] = 18'h34078; 
assign bList[153] = 18'h34306; 
assign bList[154] = 18'h34595; 
assign bList[155] = 18'h34823; 
assign bList[156] = 18'h34ab2; 
assign bList[157] = 18'h34d41; 
assign bList[158] = 18'h34fd1; 
assign bList[159] = 18'h35260; 
assign bList[160] = 18'h354ee; 
assign bList[161] = 18'h3577d; 
assign bList[162] = 18'h35a0b; 
assign bList[163] = 18'h35c98; 
assign bList[164] = 18'h35f25; 
assign bList[165] = 18'h361b1; 
assign bList[166] = 18'h3643c; 
assign bList[167] = 18'h366c6; 
assign bList[168] = 18'h3694f; 
assign bList[169] = 18'h36bd6; 
assign bList[170] = 18'h36e5c; 
assign bList[171] = 18'h370e0; 
assign bList[172] = 18'h37363; 
assign bList[173] = 18'h375e4; 
assign bList[174] = 18'h37862; 
assign bList[175] = 18'h37ade; 
assign bList[176] = 18'h37d59; 
assign bList[177] = 18'h37fd0; 
assign bList[178] = 18'h38245; 
assign bList[179] = 18'h384b7; 
assign bList[180] = 18'h38727; 
assign bList[181] = 18'h38993; 
assign bList[182] = 18'h38bfc; 
assign bList[183] = 18'h38e62; 
assign bList[184] = 18'h390c5; 
assign bList[185] = 18'h39323; 
assign bList[186] = 18'h3957e; 
assign bList[187] = 18'h397d5; 
assign bList[188] = 18'h39a28; 
assign bList[189] = 18'h39c77; 
assign bList[190] = 18'h39ec2; 
assign bList[191] = 18'h3a108; 
assign bList[192] = 18'h3a349; 
assign bList[193] = 18'h3a586; 
assign bList[194] = 18'h3a7bd; 
assign bList[195] = 18'h3a9f0; 
assign bList[196] = 18'h3ac1e; 
assign bList[197] = 18'h3ae46; 
assign bList[198] = 18'h3b068; 
assign bList[199] = 18'h3b285; 
assign bList[200] = 18'h3b49d; 
assign bList[201] = 18'h3b6ae; 
assign bList[202] = 18'h3b8ba; 
assign bList[203] = 18'h3babf; 
assign bList[204] = 18'h3bcbe; 
assign bList[205] = 18'h3beb6; 
assign bList[206] = 18'h3c0a9; 
assign bList[207] = 18'h3c294; 
assign bList[208] = 18'h3c479; 
assign bList[209] = 18'h3c657; 
assign bList[210] = 18'h3c82e; 
assign bList[211] = 18'h3c9fe; 
assign bList[212] = 18'h3cbc7; 
assign bList[213] = 18'h3cd88; 
assign bList[214] = 18'h3cf42; 
assign bList[215] = 18'h3d0f5; 
assign bList[216] = 18'h3d2a0; 
assign bList[217] = 18'h3d443; 
assign bList[218] = 18'h3d5df; 
assign bList[219] = 18'h3d773; 
assign bList[220] = 18'h3d8ff; 
assign bList[221] = 18'h3da83; 
assign bList[222] = 18'h3dc00; 
assign bList[223] = 18'h3dd74; 
assign bList[224] = 18'h3dee0; 
assign bList[225] = 18'h3e044; 
assign bList[226] = 18'h3e19f; 
assign bList[227] = 18'h3e2f3; 
assign bList[228] = 18'h3e43e; 
assign bList[229] = 18'h3e581; 
assign bList[230] = 18'h3e6bc; 
assign bList[231] = 18'h3e7ee; 
assign bList[232] = 18'h3e918; 
assign bList[233] = 18'h3ea39; 
assign bList[234] = 18'h3eb53; 
assign bList[235] = 18'h3ec64; 
assign bList[236] = 18'h3ed6c; 
assign bList[237] = 18'h3ee6d; 
assign bList[238] = 18'h3ef65; 
assign bList[239] = 18'h3f055; 
assign bList[240] = 18'h3f13c; 
assign bList[241] = 18'h3f21c; 
assign bList[242] = 18'h3f2f3; 
assign bList[243] = 18'h3f3c3; 
assign bList[244] = 18'h3f48a; 
assign bList[245] = 18'h3f54a; 
assign bList[246] = 18'h3f601; 
assign bList[247] = 18'h3f6b1; 
assign bList[248] = 18'h3f75a; 
assign bList[249] = 18'h3f7fa; 
assign bList[250] = 18'h3f894; 
assign bList[251] = 18'h3f926; 
assign bList[252] = 18'h3f9b1; 
assign bList[253] = 18'h3fa34; 
assign bList[254] = 18'h3fab1; 
assign bList[255] = 18'h3fb27; 
assign bList[256] = 18'h3fb96; 
assign bList[257] = 18'h3fbff; 
assign bList[258] = 18'h3fc61; 
assign bList[259] = 18'h3fcbd; 
assign bList[260] = 18'h3fd13; 
assign bList[261] = 18'h3fd63; 
assign bList[262] = 18'h3fdad; 
assign bList[263] = 18'h3fdf2; 
assign bList[264] = 18'h3fe31; 
assign bList[265] = 18'h3fe87; 
assign bList[266] = 18'h3fee8; 
assign bList[267] = 18'h3ff37; 
assign bList[268] = 18'h3ff76; 
assign bList[269] = 18'h3ffa6; 
assign bList[270] = 18'h3ffc9; 
assign bList[271] = 18'h3ffe2; 
assign bList[272] = 18'h3fff2; 
assign bList[273] = 18'h3fffb; 
assign bList[274] = 18'h00000; 
assign bList[275] = 18'h00000; 
assign bList[276] = 18'h00005; 
assign bList[277] = 18'h0000e; 
assign bList[278] = 18'h0001e; 
assign bList[279] = 18'h00037; 
assign bList[280] = 18'h0005a; 
assign bList[281] = 18'h0008a; 
assign bList[282] = 18'h000c9; 
assign bList[283] = 18'h00118; 
assign bList[284] = 18'h00179; 
assign bList[285] = 18'h001cf; 
assign bList[286] = 18'h0020e; 
assign bList[287] = 18'h00253; 
assign bList[288] = 18'h0029d; 
assign bList[289] = 18'h002ed; 
assign bList[290] = 18'h00343; 
assign bList[291] = 18'h0039f; 
assign bList[292] = 18'h00401; 
assign bList[293] = 18'h0046a; 
assign bList[294] = 18'h004d9; 
assign bList[295] = 18'h0054f; 
assign bList[296] = 18'h005cc; 
assign bList[297] = 18'h0064f; 
assign bList[298] = 18'h006da; 
assign bList[299] = 18'h0076c; 
assign bList[300] = 18'h00806; 
assign bList[301] = 18'h008a6; 
assign bList[302] = 18'h0094f; 
assign bList[303] = 18'h009ff; 
assign bList[304] = 18'h00ab6; 
assign bList[305] = 18'h00b76; 
assign bList[306] = 18'h00c3d; 
assign bList[307] = 18'h00d0d; 
assign bList[308] = 18'h00de4; 
assign bList[309] = 18'h00ec4; 
assign bList[310] = 18'h00fab; 
assign bList[311] = 18'h0109b; 
assign bList[312] = 18'h01193; 
assign bList[313] = 18'h01294; 
assign bList[314] = 18'h0139c; 
assign bList[315] = 18'h014ad; 
assign bList[316] = 18'h015c7; 
assign bList[317] = 18'h016e8; 
assign bList[318] = 18'h01812; 
assign bList[319] = 18'h01944; 
assign bList[320] = 18'h01a7f; 
assign bList[321] = 18'h01bc2; 
assign bList[322] = 18'h01d0d; 
assign bList[323] = 18'h01e61; 
assign bList[324] = 18'h01fbc; 
assign bList[325] = 18'h02120; 
assign bList[326] = 18'h0228c; 
assign bList[327] = 18'h02400; 
assign bList[328] = 18'h0257d; 
assign bList[329] = 18'h02701; 
assign bList[330] = 18'h0288d; 
assign bList[331] = 18'h02a21; 
assign bList[332] = 18'h02bbd; 
assign bList[333] = 18'h02d60; 
assign bList[334] = 18'h02f0b; 
assign bList[335] = 18'h030be; 
assign bList[336] = 18'h03278; 
assign bList[337] = 18'h03439; 
assign bList[338] = 18'h03602; 
assign bList[339] = 18'h037d2; 
assign bList[340] = 18'h039a9; 
assign bList[341] = 18'h03b87; 
assign bList[342] = 18'h03d6c; 
assign bList[343] = 18'h03f57; 
assign bList[344] = 18'h0414a; 
assign bList[345] = 18'h04342; 
assign bList[346] = 18'h04541; 
assign bList[347] = 18'h04746; 
assign bList[348] = 18'h04952; 
assign bList[349] = 18'h04b63; 
assign bList[350] = 18'h04d7b; 
assign bList[351] = 18'h04f98; 
assign bList[352] = 18'h051ba; 
assign bList[353] = 18'h053e2; 
assign bList[354] = 18'h05610; 
assign bList[355] = 18'h05843; 
assign bList[356] = 18'h05a7a; 
assign bList[357] = 18'h05cb7; 
assign bList[358] = 18'h05ef8; 
assign bList[359] = 18'h0613e; 
assign bList[360] = 18'h06389; 
assign bList[361] = 18'h065d8; 
assign bList[362] = 18'h0682b; 
assign bList[363] = 18'h06a82; 
assign bList[364] = 18'h06cdd; 
assign bList[365] = 18'h06f3b; 
assign bList[366] = 18'h0719e; 
assign bList[367] = 18'h07404; 
assign bList[368] = 18'h0766d; 
assign bList[369] = 18'h078d9; 
assign bList[370] = 18'h07b49; 
assign bList[371] = 18'h07dbb; 
assign bList[372] = 18'h08030; 
assign bList[373] = 18'h082a7; 
assign bList[374] = 18'h08522; 
assign bList[375] = 18'h0879e; 
assign bList[376] = 18'h08a1c; 
assign bList[377] = 18'h08c9d; 
assign bList[378] = 18'h08f20; 
assign bList[379] = 18'h091a4; 
assign bList[380] = 18'h0942a; 
assign bList[381] = 18'h096b1; 
assign bList[382] = 18'h0993a; 
assign bList[383] = 18'h09bc4; 
assign bList[384] = 18'h09e4f; 
assign bList[385] = 18'h0a0db; 
assign bList[386] = 18'h0a368; 
assign bList[387] = 18'h0a5f5; 
assign bList[388] = 18'h0a883; 
assign bList[389] = 18'h0ab12; 
assign bList[390] = 18'h0ada0; 
assign bList[391] = 18'h0b02f; 
assign bList[392] = 18'h0b2bf; 
assign bList[393] = 18'h0b54e; 
assign bList[394] = 18'h0b7dd; 
assign bList[395] = 18'h0ba6b; 
assign bList[396] = 18'h0bcfa; 
assign bList[397] = 18'h0bf88; 
assign bList[398] = 18'h0c215; 
assign bList[399] = 18'h0c4a1; 
assign bList[400] = 18'h0c72d; 
assign bList[401] = 18'h0c9b8; 
assign bList[402] = 18'h0cc42; 
assign bList[403] = 18'h0ceca; 
assign bList[404] = 18'h0d152; 
assign bList[405] = 18'h0d3d8; 
assign bList[406] = 18'h0d65d; 
assign bList[407] = 18'h0d8e0; 
assign bList[408] = 18'h0db62; 
assign bList[409] = 18'h0dde2; 
assign bList[410] = 18'h0e061; 
assign bList[411] = 18'h0e2dd; 
assign bList[412] = 18'h0e558; 
assign bList[413] = 18'h0e7d1; 
assign bList[414] = 18'h0ea47; 
assign bList[415] = 18'h0ecbc; 
assign bList[416] = 18'h0ef2e; 
assign bList[417] = 18'h0f19e; 
assign bList[418] = 18'h0f40c; 
assign bList[419] = 18'h0f677; 
assign bList[420] = 18'h0f8e0; 
assign bList[421] = 18'h0fb46; 
assign bList[422] = 18'h0fdaa; 
assign bList[423] = 18'h1000a; 
assign bList[424] = 18'h10269; 
assign bList[425] = 18'h104c4; 
assign bList[426] = 18'h1071d; 
assign bList[427] = 18'h10973; 
assign bList[428] = 18'h10bc5; 
assign bList[429] = 18'h10e15; 
assign bList[430] = 18'h11062; 
assign bList[431] = 18'h112ac; 
assign bList[432] = 18'h114f2; 
assign bList[433] = 18'h11736; 
assign bList[434] = 18'h11976; 
assign bList[435] = 18'h11bb3; 
assign bList[436] = 18'h11ded; 
assign bList[437] = 18'h12023; 
assign bList[438] = 18'h12256; 
assign bList[439] = 18'h12486; 
assign bList[440] = 18'h126b2; 
assign bList[441] = 18'h128db; 
assign bList[442] = 18'h12b00; 
assign bList[443] = 18'h12d22; 
assign bList[444] = 18'h12f41; 
assign bList[445] = 18'h1315c; 
assign bList[446] = 18'h13373; 
assign bList[447] = 18'h13587; 
assign bList[448] = 18'h13797; 
assign bList[449] = 18'h139a3; 
assign bList[450] = 18'h13bac; 
assign bList[451] = 18'h13db1; 
assign bList[452] = 18'h13fb3; 
assign bList[453] = 18'h141b1; 
assign bList[454] = 18'h143ab; 
assign bList[455] = 18'h1469a; 
assign bList[456] = 18'h14a78; 
assign bList[457] = 18'h14e47; 
assign bList[458] = 18'h15207; 
assign bList[459] = 18'h155b8; 
assign bList[460] = 18'h1595b; 
assign bList[461] = 18'h15cee; 
assign bList[462] = 18'h16072; 
assign bList[463] = 18'h163e7; 
assign bList[464] = 18'h1674e; 
assign bList[465] = 18'h16aa5; 
assign bList[466] = 18'h16dee; 
assign bList[467] = 18'h17128; 
assign bList[468] = 18'h17454; 
assign bList[469] = 18'h17770; 
assign bList[470] = 18'h17a7f; 
assign bList[471] = 18'h17d7f; 
assign bList[472] = 18'h18070; 
assign bList[473] = 18'h18354; 
assign bList[474] = 18'h1862a; 
assign bList[475] = 18'h188f2; 
assign bList[476] = 18'h18bac; 
assign bList[477] = 18'h18e59; 
assign bList[478] = 18'h190f8; 
assign bList[479] = 18'h1938a; 
assign bList[480] = 18'h1960f; 
assign bList[481] = 18'h19887; 
assign bList[482] = 18'h19af2; 
assign bList[483] = 18'h19d51; 
assign bList[484] = 18'h19fa3; 
assign bList[485] = 18'h1a1e9; 
assign bList[486] = 18'h1a423; 
assign bList[487] = 18'h1a651; 
assign bList[488] = 18'h1a873; 
assign bList[489] = 18'h1aa8a; 
assign bList[490] = 18'h1ac95; 
assign bList[491] = 18'h1ae95; 
assign bList[492] = 18'h1b08a; 
assign bList[493] = 18'h1b275; 
assign bList[494] = 18'h1b454; 
assign bList[495] = 18'h1b62a; 
assign bList[496] = 18'h1b7f4; 
assign bList[497] = 18'h1b9b5; 
assign bList[498] = 18'h1bb6c; 
assign bList[499] = 18'h1bd19; 
assign bList[500] = 18'h1bebd; 
assign bList[501] = 18'h1c057; 
assign bList[502] = 18'h1c1e8; 
assign bList[503] = 18'h1c36f; 
assign bList[504] = 18'h1c4ee; 
assign bList[505] = 18'h1c71a; 
assign bList[506] = 18'h1c9e5; 
assign bList[507] = 18'h1cc8f; 
assign bList[508] = 18'h1cf19; 
assign bList[509] = 18'h1d186; 
assign bList[510] = 18'h1d3d6; 
assign bList[511] = 18'h1d60a; 
assign bList[512] = 18'h1d823; 
assign bList[513] = 18'h1da23; 
assign bList[514] = 18'h1dc0b; 
assign bList[515] = 18'h1dddb; 
assign bList[516] = 18'h1df95; 
assign bList[517] = 18'h1e13a; 
assign bList[518] = 18'h1e2cb; 
assign bList[519] = 18'h1e448; 
assign bList[520] = 18'h1e5b2; 
assign bList[521] = 18'h1e70b; 
assign bList[522] = 18'h1e853; 
assign bList[523] = 18'h1e98a; 
assign bList[524] = 18'h1eab2; 
assign bList[525] = 18'h1ebcc; 
assign bList[526] = 18'h1ecd7; 
assign bList[527] = 18'h1edd5; 
assign bList[528] = 18'h1ef38; 
assign bList[529] = 18'h1f0ec; 
assign bList[530] = 18'h1f275; 
assign bList[531] = 18'h1f3d6; 
assign bList[532] = 18'h1f515; 
assign bList[533] = 18'h1f634; 
assign bList[534] = 18'h1f736; 
assign bList[535] = 18'h1f81e; 
assign bList[536] = 18'h1f8ef; 
assign bList[537] = 18'h1f9aa; 
assign bList[538] = 18'h1fa9d; 
assign bList[539] = 18'h1fbae; 
assign bList[540] = 18'h1fc89; 
assign bList[541] = 18'h1fd3a; 
assign bList[542] = 18'h1fdc8; 
assign bList[543] = 18'h1fe66; 
assign bList[544] = 18'h1fefb; 
assign bList[545] = 18'h1ff5a; 
assign bList[546] = 18'h1ffa9; 
assign bList[547] = 18'h1ffdd; 
assign bList[548] = 18'h1fffa; 

AND_2_1 AND_2_1_inst(
.IN_1   (   en      ),
.IN_0   (   rst_n   ),
.OUT    (   EN      )
);

always @* begin
    if(EN == 1'b1) begin
        a = aList[i];
    end
    else begin
        a = 'd0;
    end
end

always @* begin
    if(EN == 1'b1) begin
        b = bList[i];
    end
    else begin
        b = 'd0;
    end
end

endmodule
