module halfXListShift_sigmoid #(
parameter xDW = 24,
parameter ML = 196,
parameter MW = 8
)(
input wire [(MW - 1) : 0] j, //����5λ�޷�����
output wire [(xDW - 1) : 0] half_j,
output wire [(xDW - 1) : 0] half_j_1
);

wire [(xDW - 1) : 0] halfXList [(ML + 1):0]; 

// assign halfXList[0] = 16'h0000;
// assign halfXList[1] = 16'h0000;
// assign halfXList[2] = 16'h0200;
// assign halfXList[3] = 16'h0400;
// assign halfXList[4] = 16'h0600;
// assign halfXList[5] = 16'h0800;
// assign halfXList[6] = 16'h0a00;
// assign halfXList[7] = 16'h0c00;
// assign halfXList[8] = 16'h0e00;
// assign halfXList[9] = 16'h1000;
// assign halfXList[10] = 16'h1200;
// assign halfXList[11] = 16'h1400;
// assign halfXList[12] = 16'h1600;
// assign halfXList[13] = 16'h1800;
// assign halfXList[14] = 16'h1a00;
// assign halfXList[15] = 16'h1c00;
// assign halfXList[16] = 16'h2000;
// assign halfXList[17] = 16'h2400;
// assign halfXList[18] = 16'h2800;
// assign halfXList[19] = 16'h3000;
// assign halfXList[20] = 16'h4000;
// assign halfXList[21] = 16'h8000; //��Ϊ�����ʾ


// assign halfXList[0] = 24'h000000;
// assign halfXList[1] = 24'h000000; 
// assign halfXList[2] = 24'h001000; 
// assign halfXList[3] = 24'h002000; 
// assign halfXList[4] = 24'h003000; 
// assign halfXList[5] = 24'h004000; 
// assign halfXList[6] = 24'h005000; 
// assign halfXList[7] = 24'h006000; 
// assign halfXList[8] = 24'h007000; 
// assign halfXList[9] = 24'h008000; 
// assign halfXList[10] = 24'h009000; 
// assign halfXList[11] = 24'h00a000; 
// assign halfXList[12] = 24'h00b000; 
// assign halfXList[13] = 24'h00c000; 
// assign halfXList[14] = 24'h00d000; 
// assign halfXList[15] = 24'h00e000; 
// assign halfXList[16] = 24'h010000; 
// assign halfXList[17] = 24'h012000; 
// assign halfXList[18] = 24'h014000; 
// assign halfXList[19] = 24'h018000; 
// assign halfXList[20] = 24'h020000; 
// assign halfXList[21] = 24'h040000; 

assign halfXList[0] = 24'h000000; 
assign halfXList[1] = 24'h000000; 
assign halfXList[2] = 24'h000400; 
assign halfXList[3] = 24'h000800; 
assign halfXList[4] = 24'h000c00; 
assign halfXList[5] = 24'h000e00; 
assign halfXList[6] = 24'h001000; 
assign halfXList[7] = 24'h001200; 
assign halfXList[8] = 24'h001400; 
assign halfXList[9] = 24'h001600; 
assign halfXList[10] = 24'h001800; 
assign halfXList[11] = 24'h001a00; 
assign halfXList[12] = 24'h001c00; 
assign halfXList[13] = 24'h001e00; 
assign halfXList[14] = 24'h002000; 
assign halfXList[15] = 24'h002200; 
assign halfXList[16] = 24'h002400; 
assign halfXList[17] = 24'h002600; 
assign halfXList[18] = 24'h002800; 
assign halfXList[19] = 24'h002a00; 
assign halfXList[20] = 24'h002c00; 
assign halfXList[21] = 24'h002e00; 
assign halfXList[22] = 24'h003000; 
assign halfXList[23] = 24'h003200; 
assign halfXList[24] = 24'h003400; 
assign halfXList[25] = 24'h003500; 
assign halfXList[26] = 24'h003600; 
assign halfXList[27] = 24'h003700; 
assign halfXList[28] = 24'h003800; 
assign halfXList[29] = 24'h003900; 
assign halfXList[30] = 24'h003a00; 
assign halfXList[31] = 24'h003b00; 
assign halfXList[32] = 24'h003c00; 
assign halfXList[33] = 24'h003d00; 
assign halfXList[34] = 24'h003e00; 
assign halfXList[35] = 24'h003f00; 
assign halfXList[36] = 24'h004000; 
assign halfXList[37] = 24'h004100; 
assign halfXList[38] = 24'h004200; 
assign halfXList[39] = 24'h004300; 
assign halfXList[40] = 24'h004400; 
assign halfXList[41] = 24'h004500; 
assign halfXList[42] = 24'h004600; 
assign halfXList[43] = 24'h004700; 
assign halfXList[44] = 24'h004800; 
assign halfXList[45] = 24'h004900; 
assign halfXList[46] = 24'h004a00; 
assign halfXList[47] = 24'h004b00; 
assign halfXList[48] = 24'h004c00; 
assign halfXList[49] = 24'h004d00; 
assign halfXList[50] = 24'h004e00; 
assign halfXList[51] = 24'h004f00; 
assign halfXList[52] = 24'h005000; 
assign halfXList[53] = 24'h005100; 
assign halfXList[54] = 24'h005200; 
assign halfXList[55] = 24'h005300; 
assign halfXList[56] = 24'h005400; 
assign halfXList[57] = 24'h005500; 
assign halfXList[58] = 24'h005600; 
assign halfXList[59] = 24'h005700; 
assign halfXList[60] = 24'h005800; 
assign halfXList[61] = 24'h005900; 
assign halfXList[62] = 24'h005a00; 
assign halfXList[63] = 24'h005b00; 
assign halfXList[64] = 24'h005c00; 
assign halfXList[65] = 24'h005d00; 
assign halfXList[66] = 24'h005e00; 
assign halfXList[67] = 24'h005f00; 
assign halfXList[68] = 24'h006000; 
assign halfXList[69] = 24'h006100; 
assign halfXList[70] = 24'h006200; 
assign halfXList[71] = 24'h006300; 
assign halfXList[72] = 24'h006400; 
assign halfXList[73] = 24'h006500; 
assign halfXList[74] = 24'h006600; 
assign halfXList[75] = 24'h006700; 
assign halfXList[76] = 24'h006800; 
assign halfXList[77] = 24'h006900; 
assign halfXList[78] = 24'h006a00; 
assign halfXList[79] = 24'h006b00; 
assign halfXList[80] = 24'h006c00; 
assign halfXList[81] = 24'h006d00; 
assign halfXList[82] = 24'h006e00; 
assign halfXList[83] = 24'h006f00; 
assign halfXList[84] = 24'h007000; 
assign halfXList[85] = 24'h007100; 
assign halfXList[86] = 24'h007200; 
assign halfXList[87] = 24'h007300; 
assign halfXList[88] = 24'h007400; 
assign halfXList[89] = 24'h007500; 
assign halfXList[90] = 24'h007600; 
assign halfXList[91] = 24'h007700; 
assign halfXList[92] = 24'h007800; 
assign halfXList[93] = 24'h007900; 
assign halfXList[94] = 24'h007a00; 
assign halfXList[95] = 24'h007b00; 
assign halfXList[96] = 24'h007c00; 
assign halfXList[97] = 24'h007e00; 
assign halfXList[98] = 24'h008000; 
assign halfXList[99] = 24'h008200; 
assign halfXList[100] = 24'h008400; 
assign halfXList[101] = 24'h008600; 
assign halfXList[102] = 24'h008800; 
assign halfXList[103] = 24'h008a00; 
assign halfXList[104] = 24'h008c00; 
assign halfXList[105] = 24'h008e00; 
assign halfXList[106] = 24'h009000; 
assign halfXList[107] = 24'h009200; 
assign halfXList[108] = 24'h009400; 
assign halfXList[109] = 24'h009600; 
assign halfXList[110] = 24'h009800; 
assign halfXList[111] = 24'h009a00; 
assign halfXList[112] = 24'h009c00; 
assign halfXList[113] = 24'h009e00; 
assign halfXList[114] = 24'h00a000; 
assign halfXList[115] = 24'h00a200; 
assign halfXList[116] = 24'h00a400; 
assign halfXList[117] = 24'h00a600; 
assign halfXList[118] = 24'h00a800; 
assign halfXList[119] = 24'h00aa00; 
assign halfXList[120] = 24'h00ac00; 
assign halfXList[121] = 24'h00ae00; 
assign halfXList[122] = 24'h00b000; 
assign halfXList[123] = 24'h00b200; 
assign halfXList[124] = 24'h00b400; 
assign halfXList[125] = 24'h00b600; 
assign halfXList[126] = 24'h00b800; 
assign halfXList[127] = 24'h00ba00; 
assign halfXList[128] = 24'h00bc00; 
assign halfXList[129] = 24'h00be00; 
assign halfXList[130] = 24'h00c000; 
assign halfXList[131] = 24'h00c200; 
assign halfXList[132] = 24'h00c400; 
assign halfXList[133] = 24'h00c600; 
assign halfXList[134] = 24'h00c800; 
assign halfXList[135] = 24'h00ca00; 
assign halfXList[136] = 24'h00cc00; 
assign halfXList[137] = 24'h00ce00; 
assign halfXList[138] = 24'h00d000; 
assign halfXList[139] = 24'h00d200; 
assign halfXList[140] = 24'h00d400; 
assign halfXList[141] = 24'h00d600; 
assign halfXList[142] = 24'h00d800; 
assign halfXList[143] = 24'h00da00; 
assign halfXList[144] = 24'h00dc00; 
assign halfXList[145] = 24'h00de00; 
assign halfXList[146] = 24'h00e000; 
assign halfXList[147] = 24'h00e200; 
assign halfXList[148] = 24'h00e400; 
assign halfXList[149] = 24'h00e600; 
assign halfXList[150] = 24'h00e800; 
assign halfXList[151] = 24'h00ea00; 
assign halfXList[152] = 24'h00ec00; 
assign halfXList[153] = 24'h00ee00; 
assign halfXList[154] = 24'h00f000; 
assign halfXList[155] = 24'h00f200; 
assign halfXList[156] = 24'h00f400; 
assign halfXList[157] = 24'h00f800; 
assign halfXList[158] = 24'h00fc00; 
assign halfXList[159] = 24'h010000; 
assign halfXList[160] = 24'h010400; 
assign halfXList[161] = 24'h010800; 
assign halfXList[162] = 24'h010c00; 
assign halfXList[163] = 24'h011000; 
assign halfXList[164] = 24'h011400; 
assign halfXList[165] = 24'h011800; 
assign halfXList[166] = 24'h011c00; 
assign halfXList[167] = 24'h012000; 
assign halfXList[168] = 24'h012400; 
assign halfXList[169] = 24'h012800; 
assign halfXList[170] = 24'h012c00; 
assign halfXList[171] = 24'h013000; 
assign halfXList[172] = 24'h013400; 
assign halfXList[173] = 24'h013800; 
assign halfXList[174] = 24'h013c00; 
assign halfXList[175] = 24'h014000; 
assign halfXList[176] = 24'h014400; 
assign halfXList[177] = 24'h014800; 
assign halfXList[178] = 24'h014c00; 
assign halfXList[179] = 24'h015000; 
assign halfXList[180] = 24'h015800; 
assign halfXList[181] = 24'h016000; 
assign halfXList[182] = 24'h016800; 
assign halfXList[183] = 24'h017000; 
assign halfXList[184] = 24'h017800; 
assign halfXList[185] = 24'h018000; 
assign halfXList[186] = 24'h018800; 
assign halfXList[187] = 24'h019000; 
assign halfXList[188] = 24'h019800; 
assign halfXList[189] = 24'h01a000; 
assign halfXList[190] = 24'h01a800; 
assign halfXList[191] = 24'h01b000; 
assign halfXList[192] = 24'h01c000; 
assign halfXList[193] = 24'h01d000; 
assign halfXList[194] = 24'h01e000; 
assign halfXList[195] = 24'h01f000; 
assign halfXList[196] = 24'h020000; 
assign halfXList[197] = 24'h040000;

assign half_j = halfXList[j];
assign half_j_1 = halfXList[j + 1'b1];

endmodule