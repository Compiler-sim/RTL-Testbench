module wi_buffer #(
  parameter D_WL = 24,
  parameter UNITS_NUM = 5
)(
   input [7:0] addr,
   output [UNITS_NUM*D_WL-1:0] w_o
);

wire [D_WL*UNITS_NUM-1:0] w_fix [0:155];
assign w_o = w_fix[addr];
assign w_fix[0]='hffff57000846ffffe9fffef00003a4;
assign w_fix[1]='hfff78e000809fff75efff345000807;
assign w_fix[2]='hffece1001ff9ffefeeffed7ffffa97;
assign w_fix[3]='hffef280004d3ffd585ffebeaffefd5;
assign w_fix[4]='hfff201ffde3afff665fff5ceffd2e6;
assign w_fix[5]='hffe8e1000568ffeb78fff3f0fff732;
assign w_fix[6]='hffeaef000f57fffeb7fffd47002108;
assign w_fix[7]='hfffd970024ec0000b7fff890003fac;
assign w_fix[8]='hfffb920004c6fff073fff369003321;
assign w_fix[9]='h00013c000429ffea5ffff1eb002fc3;
assign w_fix[10]='h00002e001aa100031400038a000e54;
assign w_fix[11]='hfffbd1fffa5bfffff6fffdc5001e74;
assign w_fix[12]='hfffe2efff6120000f6fffbd800127d;
assign w_fix[13]='hfffb3afffa23fffb13fffacf0011ec;
assign w_fix[14]='hfffbf6fffeb0fffbaffff6d4001dbf;
assign w_fix[15]='hfffc6efffad80015e8ffedf0002cf0;
assign w_fix[16]='hfffd0fffe7f0002050ffebde001edb;
assign w_fix[17]='hfffa0bffe6b70013c6fff190002240;
assign w_fix[18]='hfff84bffbc01000d3fffead1003320;
assign w_fix[19]='hfffd06ffe153000795fff243004182;
assign w_fix[20]='hfffb170005cafff8e7fff201004fe5;
assign w_fix[21]='hfff68d000e55ffe9d1fff593003596;
assign w_fix[22]='hfff2f5000f1ffff627fff881001d8e;
assign w_fix[23]='hffeeff00065fffed84fff9a2002040;
assign w_fix[24]='hfff6a50002b6ffee65fff7f20027e2;
assign w_fix[25]='hfffa93fffac7fff82efffb82000897;
assign w_fix[26]='hfffee1fffa80000012ffef160002ac;
assign w_fix[27]='hfff151ffefe3fffe35ffde96000220;
assign w_fix[28]='hfffb42ffce00fff46fffe9d2000b0c;
assign w_fix[29]='hffdd44ffe11ffff7adffe7ec000c2f;
assign w_fix[30]='h0011ccfff228ffffba0004950010e1;
assign w_fix[31]='hfff6390019c300055afff617000a1f;
assign w_fix[32]='hfff20d001a6c000cefffe1c7000623;
assign w_fix[33]='hfff0a0000e21fffb61ffd6cffff711;
assign w_fix[34]='hfff1a9001a5afff9dbffe4aefffe81;
assign w_fix[35]='hffe8630015f0fffa62fff72300040d;
assign w_fix[36]='h0001cd000f570006b3fff3ed000460;
assign w_fix[37]='hfffb78000f27ffff51ffe75afff920;
assign w_fix[38]='hfffeb7000c8400026affdf16fff58f;
assign w_fix[39]='h000598fffbe10004ccffdefdffecec;
assign w_fix[40]='hffff1afffc2500022bffe2aaffef51;
assign w_fix[41]='h00132cfffcd70001cdffdbbcffec36;
assign w_fix[42]='h001d59fff8b300007dffe34affed0c;
assign w_fix[43]='h001a6a000aa000091bffe359fff7cc;
assign w_fix[44]='hfffb9ffff0f2000b2efff589fff3a1;
assign w_fix[45]='hffffa4ffee4f000831000297fffff0;
assign w_fix[46]='hfffea7fff9f6000d59fffb7d000f16;
assign w_fix[47]='hfff72d00059b000a28ffe186000958;
assign w_fix[48]='h000012001253000633ffe480fff962;
assign w_fix[49]='h00083400186afff9adffe83bfff320;
assign w_fix[50]='h000926fff54ffff3d8fff06300023f;
assign w_fix[51]='hffffedffe6fdfffb22ffebc4000176;
assign w_fix[52]='h000004fffd3dffff53000838000004;
assign w_fix[53]='hfffff5fff532fff07e001570ffffc4;
assign w_fix[54]='hfffffaffe853fff383000148fffbcf;
assign w_fix[55]='hffff6afff4c6ffe6e2003616fffa5f;
assign w_fix[56]='hfffedbfff687001445fffe68fffb64;
assign w_fix[57]='hffff3a0014a3fff806002f4bfff7d0;
assign w_fix[58]='hfffd2a000f74fff0170016befffafa;
assign w_fix[59]='hffff85fffb5fffec80fffdf9fff8c9;
assign w_fix[60]='hfffe280000c4fff267ffff92fffa32;
assign w_fix[61]='hfffdcc00092afff7e90012d7fffb69;
assign w_fix[62]='hffff50000527001bd200008ffffdf1;
assign w_fix[63]='hffffd6fffbdffff72300096cfffdb8;
assign w_fix[64]='hffffd8000bd9ffff53001173fffd8a;
assign w_fix[65]='hffff78000028000918000a9dfffecf;
assign w_fix[66]='hffff83fffbe8ffff5b0008f4ffff70;
assign w_fix[67]='hfffed8fff67a0009bbfff3f1fffdb2;
assign w_fix[68]='hfffd9cfff142000779ffe27efffb41;
assign w_fix[69]='hfffe140004660012c5ffe2defffaf7;
assign w_fix[70]='hfffd21002397fff73dffeb22fff97f;
assign w_fix[71]='hfffeda002d010004e9ffecc5fffd6e;
assign w_fix[72]='hfffe0f0011d300144cfff555fffc51;
assign w_fix[73]='hfffd3d001881000bcc0003cafffd33;
assign w_fix[74]='hfffd2b0016ef000e52001233fffe96;
assign w_fix[75]='hfffc910009c000088f000820ffff49;
assign w_fix[76]='hfffd93000b53000776001067fffe99;
assign w_fix[77]='hffff27000a82ffffb3001e45fffff0;
assign w_fix[78]='h00004b0000fcffff96fff93fffeeab;
assign w_fix[79]='h00024f000612fffd9ffff45dffdbce;
assign w_fix[80]='h0004e40007c0fffe93ffe3c4ffe109;
assign w_fix[81]='h000a52000735000612ffd289ffe3ea;
assign w_fix[82]='h00065400124d000228fff4e6000022;
assign w_fix[83]='h000033001108000e02ffe286000ec7;
assign w_fix[84]='h000b7c00086000019effff840003f6;
assign w_fix[85]='h001018001367000587ffff4cffdc27;
assign w_fix[86]='h000112000b74000401000231ffec89;
assign w_fix[87]='hfffd1f0012cf00028affea530002f3;
assign w_fix[88]='h0009b100022a000391000cd8fff48e;
assign w_fix[89]='h0006840002df000549001addfff048;
assign w_fix[90]='h000278fffe49000346000ee7ffece2;
assign w_fix[91]='h0000defffded000056001996ffdfb9;
assign w_fix[92]='h00015efff1840000e1001087ffdccf;
assign w_fix[93]='h00020bffe8d2ffffd5001f12ffe1bf;
assign w_fix[94]='hfffe4d0006f90000e6001318fff83d;
assign w_fix[95]='hffff630006f2000423000714fffa91;
assign w_fix[96]='hfffd2bfff28a000414ffe0c8fffbe4;
assign w_fix[97]='h000854fff50f000618ffec890008ed;
assign w_fix[98]='h000693fff39d000535ffeff700072d;
assign w_fix[99]='h0004bcfff465000550fff7bfffdb6e;
assign w_fix[100]='h0003ddfff6c0000586fffe6dffd55e;
assign w_fix[101]='h000451fff88c0005c1000e36ffdd20;
assign w_fix[102]='h000444fff941000752fffed0ffe282;
assign w_fix[103]='h0000c2fffa9f00050fffefd8ffdf0b;
assign w_fix[104]='h000030fffd6bffe97300007afffefb;
assign w_fix[105]='hfffd70ffeb39ffe73c00027f000084;
assign w_fix[106]='h000502ffea88fff92c000a620003f0;
assign w_fix[107]='h000a49ffd61cfffab000076f00057f;
assign w_fix[108]='h00098d002af2ffee310005f9000a17;
assign w_fix[109]='h00049d0009f10003ce000733000ef5;
assign w_fix[110]='h000bb6fff5ed001e380005ba000891;
assign w_fix[111]='h0016a2ffe011000c580004f5000e49;
assign w_fix[112]='h000c29fff62cffe10f0008000013bb;
assign w_fix[113]='h0000560004120005a10001a0000f3c;
assign w_fix[114]='hfffea3001dd60007200001500009a2;
assign w_fix[115]='h0002a3fff748fff253fffffb00099a;
assign w_fix[116]='h000449fffb18fffa2ffffeba000750;
assign w_fix[117]='h0002060008260004d4ffff81fffe98;
assign w_fix[118]='h0000b5fffb74001381ffffdbfffe1a;
assign w_fix[119]='h0000cbfff9c8000c26ffff8300092b;
assign w_fix[120]='h0005e2fffe9d000aef00010b0010c5;
assign w_fix[121]='h00082ffffe4c000c45000712000678;
assign w_fix[122]='h00145bfffeb6fff16600048d000e54;
assign w_fix[123]='h0012f9000ad70009a900000a000e2e;
assign w_fix[124]='h00065f00102efff1f5fff56d000b06;
assign w_fix[125]='h000447000780ffd9a0fffee1000679;
assign w_fix[126]='h000080000e46ffee0ffffcfc000b4b;
assign w_fix[127]='h000613000e9efff9e8fffc13000776;
assign w_fix[128]='h000354000ac90008cbfffc900009cf;
assign w_fix[129]='h00038a000696ffe781fffadf000319;
assign w_fix[130]='h000009fffe1c00068efffe6afffde4;
assign w_fix[131]='h00003cfff298001a7cfff1a4ffea06;
assign w_fix[132]='hfffe24fff1c30019fbffe9a3ffe36c;
assign w_fix[133]='hfffe66ffdc240001b6fff0eaffe5a9;
assign w_fix[134]='hfffcaa00147d000dc100095cffeee5;
assign w_fix[135]='hfffc5a0005af0019c6001c18ffeaa3;
assign w_fix[136]='hfffd28ffe9beffedaf001cf3fff586;
assign w_fix[137]='hfffb3affe5f2fff302000892ffecac;
assign w_fix[138]='hfffb28fff739fffbfa0006a9fff096;
assign w_fix[139]='hfffe12fffa4d001147000b4afff310;
assign w_fix[140]='hffff1f000950ffd912000ff6ffff2a;
assign w_fix[141]='hffffeafff5c2ffcf5900072cfff823;
assign w_fix[142]='hffff7afffc57ffeaf60001e7fffa56;
assign w_fix[143]='h00003c0006a9fff97ffffe8afff334;
assign w_fix[144]='h000004ffff6bfff284fffc55fff2aa;
assign w_fix[145]='hffffea0003b9ffe90400024bffe8d7;
assign w_fix[146]='hffffe8000401ffec0d00098affe3b6;
assign w_fix[147]='h000044fff88d0000cf000ecbffe916;
assign w_fix[148]='hfffba90008b7fff6d9ffff7effe9b6;
assign w_fix[149]='hfffc6a000b90000f5bfffde4ffefe6;
assign w_fix[150]='hfffd1f0005fb0005f1fffea4fff0aa;
assign w_fix[151]='hfffe72fffe99001556fff1d2fff015;
assign w_fix[152]='hffff180004c10008ffffecc2fff238;
assign w_fix[153]='hfffee40007800021c0fffc6affed30;
assign w_fix[154]='hfffe23000773001623fffb2fffe774;
assign w_fix[155]='hffffc200040a00000ffff09cffea9c;

endmodule